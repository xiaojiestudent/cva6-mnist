//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2018/08/07 15:45:30
// Design Name: 
// Module Name: rom_pxc
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module rom_pxc(
   input clk,
   input ena,
   input [13 : 0] addr,
   output [9 : 0] dout
    );
    
    reg [9 : 0]pxcRom[0 : 15679];
    /*
    initial
    begin
       $readmemb( "C:/Users/Dell/Desktop/bayes_test_reg/p_xi_c_b.dat", pxcRom);
    end
    */
    
    always@( posedge clk)
    begin
    pxcRom[0] <= 10'b0000000000;
    pxcRom[1] <= 10'b0000000000;
    pxcRom[2] <= 10'b0000000000;
    pxcRom[3] <= 10'b0000000000;
    pxcRom[4] <= 10'b0000000000;
    pxcRom[5] <= 10'b0000000000;
    pxcRom[6] <= 10'b0000000000;
    pxcRom[7] <= 10'b0000000000;
    pxcRom[8] <= 10'b0000000000;
    pxcRom[9] <= 10'b0000000000;
    pxcRom[10] <= 10'b0000000000;
    pxcRom[11] <= 10'b0000000000;
    pxcRom[12] <= 10'b0000000000;
    pxcRom[13] <= 10'b0000000000;
    pxcRom[14] <= 10'b0000000000;
    pxcRom[15] <= 10'b0000000000;
    pxcRom[16] <= 10'b0000000000;
    pxcRom[17] <= 10'b0000000000;
    pxcRom[18] <= 10'b0000000000;
    pxcRom[19] <= 10'b0000000000;
    pxcRom[20] <= 10'b0000000000;
    pxcRom[21] <= 10'b0000000000;
    pxcRom[22] <= 10'b0000000000;
    pxcRom[23] <= 10'b0000000000;
    pxcRom[24] <= 10'b0000000000;
    pxcRom[25] <= 10'b0000000000;
    pxcRom[26] <= 10'b0000000000;
    pxcRom[27] <= 10'b0000000000;
    pxcRom[28] <= 10'b0000000000;
    pxcRom[29] <= 10'b0000000000;
    pxcRom[30] <= 10'b0000000000;
    pxcRom[31] <= 10'b0000000000;
    pxcRom[32] <= 10'b0000000000;
    pxcRom[33] <= 10'b0000000000;
    pxcRom[34] <= 10'b0000000000;
    pxcRom[35] <= 10'b0000000000;
    pxcRom[36] <= 10'b0000000000;
    pxcRom[37] <= 10'b0000000000;
    pxcRom[38] <= 10'b0000000000;
    pxcRom[39] <= 10'b0000000000;
    pxcRom[40] <= 10'b0000000000;
    pxcRom[41] <= 10'b0000000000;
    pxcRom[42] <= 10'b0000000000;
    pxcRom[43] <= 10'b0000000000;
    pxcRom[44] <= 10'b0000000000;
    pxcRom[45] <= 10'b0000000000;
    pxcRom[46] <= 10'b0000000000;
    pxcRom[47] <= 10'b0000000000;
    pxcRom[48] <= 10'b0000000000;
    pxcRom[49] <= 10'b0000000000;
    pxcRom[50] <= 10'b0000000000;
    pxcRom[51] <= 10'b0000000000;
    pxcRom[52] <= 10'b0000000000;
    pxcRom[53] <= 10'b0000000000;
    pxcRom[54] <= 10'b0000000000;
    pxcRom[55] <= 10'b0000000000;
    pxcRom[56] <= 10'b0000000000;
    pxcRom[57] <= 10'b0000000000;
    pxcRom[58] <= 10'b0000000000;
    pxcRom[59] <= 10'b0000000000;
    pxcRom[60] <= 10'b0000000000;
    pxcRom[61] <= 10'b0000000000;
    pxcRom[62] <= 10'b0000000000;
    pxcRom[63] <= 10'b0000000000;
    pxcRom[64] <= 10'b0000000000;
    pxcRom[65] <= 10'b0000000000;
    pxcRom[66] <= 10'b0000000000;
    pxcRom[67] <= 10'b0000000000;
    pxcRom[68] <= 10'b0000000000;
    pxcRom[69] <= 10'b0000000000;
    pxcRom[70] <= 10'b0000000000;
    pxcRom[71] <= 10'b0000000000;
    pxcRom[72] <= 10'b0000000000;
    pxcRom[73] <= 10'b0000000000;
    pxcRom[74] <= 10'b0000000000;
    pxcRom[75] <= 10'b0000000000;
    pxcRom[76] <= 10'b0000000000;
    pxcRom[77] <= 10'b0000000000;
    pxcRom[78] <= 10'b0000000000;
    pxcRom[79] <= 10'b0000000000;
    pxcRom[80] <= 10'b0000000000;
    pxcRom[81] <= 10'b0000000000;
    pxcRom[82] <= 10'b0000000000;
    pxcRom[83] <= 10'b0000000000;
    pxcRom[84] <= 10'b0000000000;
    pxcRom[85] <= 10'b0000000000;
    pxcRom[86] <= 10'b0000000000;
    pxcRom[87] <= 10'b0000000000;
    pxcRom[88] <= 10'b0000000000;
    pxcRom[89] <= 10'b0000000000;
    pxcRom[90] <= 10'b0000000000;
    pxcRom[91] <= 10'b0000000000;
    pxcRom[92] <= 10'b0000000000;
    pxcRom[93] <= 10'b0000000000;
    pxcRom[94] <= 10'b0000000000;
    pxcRom[95] <= 10'b0000000000;
    pxcRom[96] <= 10'b0000000000;
    pxcRom[97] <= 10'b0000000001;
    pxcRom[98] <= 10'b0000000001;
    pxcRom[99] <= 10'b0000000001;
    pxcRom[100] <= 10'b0000000001;
    pxcRom[101] <= 10'b0000000001;
    pxcRom[102] <= 10'b0000000001;
    pxcRom[103] <= 10'b0000000000;
    pxcRom[104] <= 10'b0000000000;
    pxcRom[105] <= 10'b0000000000;
    pxcRom[106] <= 10'b0000000000;
    pxcRom[107] <= 10'b0000000000;
    pxcRom[108] <= 10'b0000000000;
    pxcRom[109] <= 10'b0000000000;
    pxcRom[110] <= 10'b0000000000;
    pxcRom[111] <= 10'b0000000000;
    pxcRom[112] <= 10'b0000000000;
    pxcRom[113] <= 10'b0000000000;
    pxcRom[114] <= 10'b0000000000;
    pxcRom[115] <= 10'b0000000000;
    pxcRom[116] <= 10'b0000000000;
    pxcRom[117] <= 10'b0000000000;
    pxcRom[118] <= 10'b0000000000;
    pxcRom[119] <= 10'b0000000000;
    pxcRom[120] <= 10'b0000000000;
    pxcRom[121] <= 10'b0000000001;
    pxcRom[122] <= 10'b0000000011;
    pxcRom[123] <= 10'b0000000110;
    pxcRom[124] <= 10'b0000001011;
    pxcRom[125] <= 10'b0000010001;
    pxcRom[126] <= 10'b0000010111;
    pxcRom[127] <= 10'b0000011100;
    pxcRom[128] <= 10'b0000011101;
    pxcRom[129] <= 10'b0000011011;
    pxcRom[130] <= 10'b0000010101;
    pxcRom[131] <= 10'b0000001111;
    pxcRom[132] <= 10'b0000001001;
    pxcRom[133] <= 10'b0000000100;
    pxcRom[134] <= 10'b0000000010;
    pxcRom[135] <= 10'b0000000000;
    pxcRom[136] <= 10'b0000000000;
    pxcRom[137] <= 10'b0000000000;
    pxcRom[138] <= 10'b0000000000;
    pxcRom[139] <= 10'b0000000000;
    pxcRom[140] <= 10'b0000000000;
    pxcRom[141] <= 10'b0000000000;
    pxcRom[142] <= 10'b0000000000;
    pxcRom[143] <= 10'b0000000000;
    pxcRom[144] <= 10'b0000000000;
    pxcRom[145] <= 10'b0000000000;
    pxcRom[146] <= 10'b0000000000;
    pxcRom[147] <= 10'b0000000000;
    pxcRom[148] <= 10'b0000000010;
    pxcRom[149] <= 10'b0000000101;
    pxcRom[150] <= 10'b0000001010;
    pxcRom[151] <= 10'b0000010010;
    pxcRom[152] <= 10'b0000011111;
    pxcRom[153] <= 10'b0000101111;
    pxcRom[154] <= 10'b0000111111;
    pxcRom[155] <= 10'b0001001110;
    pxcRom[156] <= 10'b0001010011;
    pxcRom[157] <= 10'b0001001100;
    pxcRom[158] <= 10'b0000111010;
    pxcRom[159] <= 10'b0000101000;
    pxcRom[160] <= 10'b0000011001;
    pxcRom[161] <= 10'b0000001101;
    pxcRom[162] <= 10'b0000000101;
    pxcRom[163] <= 10'b0000000001;
    pxcRom[164] <= 10'b0000000000;
    pxcRom[165] <= 10'b0000000000;
    pxcRom[166] <= 10'b0000000000;
    pxcRom[167] <= 10'b0000000000;
    pxcRom[168] <= 10'b0000000000;
    pxcRom[169] <= 10'b0000000000;
    pxcRom[170] <= 10'b0000000000;
    pxcRom[171] <= 10'b0000000000;
    pxcRom[172] <= 10'b0000000000;
    pxcRom[173] <= 10'b0000000000;
    pxcRom[174] <= 10'b0000000000;
    pxcRom[175] <= 10'b0000000010;
    pxcRom[176] <= 10'b0000000101;
    pxcRom[177] <= 10'b0000001010;
    pxcRom[178] <= 10'b0000010101;
    pxcRom[179] <= 10'b0000100100;
    pxcRom[180] <= 10'b0000111000;
    pxcRom[181] <= 10'b0001010000;
    pxcRom[182] <= 10'b0001100110;
    pxcRom[183] <= 10'b0001111010;
    pxcRom[184] <= 10'b0010000001;
    pxcRom[185] <= 10'b0001111010;
    pxcRom[186] <= 10'b0001100110;
    pxcRom[187] <= 10'b0001001000;
    pxcRom[188] <= 10'b0000101101;
    pxcRom[189] <= 10'b0000011011;
    pxcRom[190] <= 10'b0000001100;
    pxcRom[191] <= 10'b0000000100;
    pxcRom[192] <= 10'b0000000000;
    pxcRom[193] <= 10'b0000000000;
    pxcRom[194] <= 10'b0000000000;
    pxcRom[195] <= 10'b0000000000;
    pxcRom[196] <= 10'b0000000000;
    pxcRom[197] <= 10'b0000000000;
    pxcRom[198] <= 10'b0000000000;
    pxcRom[199] <= 10'b0000000000;
    pxcRom[200] <= 10'b0000000000;
    pxcRom[201] <= 10'b0000000000;
    pxcRom[202] <= 10'b0000000001;
    pxcRom[203] <= 10'b0000000100;
    pxcRom[204] <= 10'b0000001010;
    pxcRom[205] <= 10'b0000010100;
    pxcRom[206] <= 10'b0000100101;
    pxcRom[207] <= 10'b0000111011;
    pxcRom[208] <= 10'b0001010011;
    pxcRom[209] <= 10'b0001101001;
    pxcRom[210] <= 10'b0001110110;
    pxcRom[211] <= 10'b0001111010;
    pxcRom[212] <= 10'b0001111111;
    pxcRom[213] <= 10'b0010000011;
    pxcRom[214] <= 10'b0001111101;
    pxcRom[215] <= 10'b0001100111;
    pxcRom[216] <= 10'b0001001000;
    pxcRom[217] <= 10'b0000101011;
    pxcRom[218] <= 10'b0000010110;
    pxcRom[219] <= 10'b0000001001;
    pxcRom[220] <= 10'b0000000001;
    pxcRom[221] <= 10'b0000000000;
    pxcRom[222] <= 10'b0000000000;
    pxcRom[223] <= 10'b0000000000;
    pxcRom[224] <= 10'b0000000000;
    pxcRom[225] <= 10'b0000000000;
    pxcRom[226] <= 10'b0000000000;
    pxcRom[227] <= 10'b0000000000;
    pxcRom[228] <= 10'b0000000000;
    pxcRom[229] <= 10'b0000000000;
    pxcRom[230] <= 10'b0000000011;
    pxcRom[231] <= 10'b0000001000;
    pxcRom[232] <= 10'b0000010010;
    pxcRom[233] <= 10'b0000100010;
    pxcRom[234] <= 10'b0000111001;
    pxcRom[235] <= 10'b0001010001;
    pxcRom[236] <= 10'b0001100011;
    pxcRom[237] <= 10'b0001100101;
    pxcRom[238] <= 10'b0001011110;
    pxcRom[239] <= 10'b0001010110;
    pxcRom[240] <= 10'b0001010011;
    pxcRom[241] <= 10'b0001011010;
    pxcRom[242] <= 10'b0001100110;
    pxcRom[243] <= 10'b0001101100;
    pxcRom[244] <= 10'b0001011011;
    pxcRom[245] <= 10'b0000111110;
    pxcRom[246] <= 10'b0000100001;
    pxcRom[247] <= 10'b0000001111;
    pxcRom[248] <= 10'b0000000011;
    pxcRom[249] <= 10'b0000000000;
    pxcRom[250] <= 10'b0000000000;
    pxcRom[251] <= 10'b0000000000;
    pxcRom[252] <= 10'b0000000000;
    pxcRom[253] <= 10'b0000000000;
    pxcRom[254] <= 10'b0000000000;
    pxcRom[255] <= 10'b0000000000;
    pxcRom[256] <= 10'b0000000000;
    pxcRom[257] <= 10'b0000000001;
    pxcRom[258] <= 10'b0000000101;
    pxcRom[259] <= 10'b0000001111;
    pxcRom[260] <= 10'b0000011101;
    pxcRom[261] <= 10'b0000110100;
    pxcRom[262] <= 10'b0001001100;
    pxcRom[263] <= 10'b0001011111;
    pxcRom[264] <= 10'b0001011110;
    pxcRom[265] <= 10'b0001001111;
    pxcRom[266] <= 10'b0000111110;
    pxcRom[267] <= 10'b0000110011;
    pxcRom[268] <= 10'b0000110000;
    pxcRom[269] <= 10'b0000110011;
    pxcRom[270] <= 10'b0001000010;
    pxcRom[271] <= 10'b0001010111;
    pxcRom[272] <= 10'b0001100010;
    pxcRom[273] <= 10'b0001001110;
    pxcRom[274] <= 10'b0000101110;
    pxcRom[275] <= 10'b0000010110;
    pxcRom[276] <= 10'b0000000101;
    pxcRom[277] <= 10'b0000000000;
    pxcRom[278] <= 10'b0000000000;
    pxcRom[279] <= 10'b0000000000;
    pxcRom[280] <= 10'b0000000000;
    pxcRom[281] <= 10'b0000000000;
    pxcRom[282] <= 10'b0000000000;
    pxcRom[283] <= 10'b0000000000;
    pxcRom[284] <= 10'b0000000000;
    pxcRom[285] <= 10'b0000000011;
    pxcRom[286] <= 10'b0000001010;
    pxcRom[287] <= 10'b0000010111;
    pxcRom[288] <= 10'b0000101100;
    pxcRom[289] <= 10'b0001000111;
    pxcRom[290] <= 10'b0001011101;
    pxcRom[291] <= 10'b0001011110;
    pxcRom[292] <= 10'b0001001010;
    pxcRom[293] <= 10'b0000110101;
    pxcRom[294] <= 10'b0000100110;
    pxcRom[295] <= 10'b0000011100;
    pxcRom[296] <= 10'b0000010111;
    pxcRom[297] <= 10'b0000011011;
    pxcRom[298] <= 10'b0000101001;
    pxcRom[299] <= 10'b0001000010;
    pxcRom[300] <= 10'b0001011011;
    pxcRom[301] <= 10'b0001011000;
    pxcRom[302] <= 10'b0000111010;
    pxcRom[303] <= 10'b0000011101;
    pxcRom[304] <= 10'b0000000111;
    pxcRom[305] <= 10'b0000000000;
    pxcRom[306] <= 10'b0000000000;
    pxcRom[307] <= 10'b0000000000;
    pxcRom[308] <= 10'b0000000000;
    pxcRom[309] <= 10'b0000000000;
    pxcRom[310] <= 10'b0000000000;
    pxcRom[311] <= 10'b0000000000;
    pxcRom[312] <= 10'b0000000000;
    pxcRom[313] <= 10'b0000000110;
    pxcRom[314] <= 10'b0000010000;
    pxcRom[315] <= 10'b0000100011;
    pxcRom[316] <= 10'b0000111101;
    pxcRom[317] <= 10'b0001011001;
    pxcRom[318] <= 10'b0001100000;
    pxcRom[319] <= 10'b0001001100;
    pxcRom[320] <= 10'b0000110100;
    pxcRom[321] <= 10'b0000100001;
    pxcRom[322] <= 10'b0000010100;
    pxcRom[323] <= 10'b0000001101;
    pxcRom[324] <= 10'b0000001011;
    pxcRom[325] <= 10'b0000001111;
    pxcRom[326] <= 10'b0000011011;
    pxcRom[327] <= 10'b0000110011;
    pxcRom[328] <= 10'b0001010001;
    pxcRom[329] <= 10'b0001011110;
    pxcRom[330] <= 10'b0001000010;
    pxcRom[331] <= 10'b0000100011;
    pxcRom[332] <= 10'b0000001010;
    pxcRom[333] <= 10'b0000000000;
    pxcRom[334] <= 10'b0000000000;
    pxcRom[335] <= 10'b0000000000;
    pxcRom[336] <= 10'b0000000000;
    pxcRom[337] <= 10'b0000000000;
    pxcRom[338] <= 10'b0000000000;
    pxcRom[339] <= 10'b0000000000;
    pxcRom[340] <= 10'b0000000001;
    pxcRom[341] <= 10'b0000001001;
    pxcRom[342] <= 10'b0000011001;
    pxcRom[343] <= 10'b0000110001;
    pxcRom[344] <= 10'b0001001111;
    pxcRom[345] <= 10'b0001100001;
    pxcRom[346] <= 10'b0001010100;
    pxcRom[347] <= 10'b0000111000;
    pxcRom[348] <= 10'b0000100001;
    pxcRom[349] <= 10'b0000010010;
    pxcRom[350] <= 10'b0000001001;
    pxcRom[351] <= 10'b0000000110;
    pxcRom[352] <= 10'b0000000101;
    pxcRom[353] <= 10'b0000001010;
    pxcRom[354] <= 10'b0000010101;
    pxcRom[355] <= 10'b0000101011;
    pxcRom[356] <= 10'b0001001011;
    pxcRom[357] <= 10'b0001011100;
    pxcRom[358] <= 10'b0001000110;
    pxcRom[359] <= 10'b0000100111;
    pxcRom[360] <= 10'b0000001100;
    pxcRom[361] <= 10'b0000000000;
    pxcRom[362] <= 10'b0000000000;
    pxcRom[363] <= 10'b0000000000;
    pxcRom[364] <= 10'b0000000000;
    pxcRom[365] <= 10'b0000000000;
    pxcRom[366] <= 10'b0000000000;
    pxcRom[367] <= 10'b0000000000;
    pxcRom[368] <= 10'b0000000010;
    pxcRom[369] <= 10'b0000001111;
    pxcRom[370] <= 10'b0000100011;
    pxcRom[371] <= 10'b0001000000;
    pxcRom[372] <= 10'b0001011101;
    pxcRom[373] <= 10'b0001011110;
    pxcRom[374] <= 10'b0001000010;
    pxcRom[375] <= 10'b0000100110;
    pxcRom[376] <= 10'b0000010011;
    pxcRom[377] <= 10'b0000001000;
    pxcRom[378] <= 10'b0000000100;
    pxcRom[379] <= 10'b0000000010;
    pxcRom[380] <= 10'b0000000011;
    pxcRom[381] <= 10'b0000001000;
    pxcRom[382] <= 10'b0000010100;
    pxcRom[383] <= 10'b0000101001;
    pxcRom[384] <= 10'b0001001000;
    pxcRom[385] <= 10'b0001011011;
    pxcRom[386] <= 10'b0001000101;
    pxcRom[387] <= 10'b0000100110;
    pxcRom[388] <= 10'b0000001100;
    pxcRom[389] <= 10'b0000000000;
    pxcRom[390] <= 10'b0000000000;
    pxcRom[391] <= 10'b0000000000;
    pxcRom[392] <= 10'b0000000000;
    pxcRom[393] <= 10'b0000000000;
    pxcRom[394] <= 10'b0000000000;
    pxcRom[395] <= 10'b0000000000;
    pxcRom[396] <= 10'b0000000011;
    pxcRom[397] <= 10'b0000010101;
    pxcRom[398] <= 10'b0000101110;
    pxcRom[399] <= 10'b0001010000;
    pxcRom[400] <= 10'b0001100100;
    pxcRom[401] <= 10'b0001010001;
    pxcRom[402] <= 10'b0000110010;
    pxcRom[403] <= 10'b0000011000;
    pxcRom[404] <= 10'b0000001010;
    pxcRom[405] <= 10'b0000000100;
    pxcRom[406] <= 10'b0000000010;
    pxcRom[407] <= 10'b0000000001;
    pxcRom[408] <= 10'b0000000011;
    pxcRom[409] <= 10'b0000001001;
    pxcRom[410] <= 10'b0000010110;
    pxcRom[411] <= 10'b0000101101;
    pxcRom[412] <= 10'b0001001010;
    pxcRom[413] <= 10'b0001010111;
    pxcRom[414] <= 10'b0001000000;
    pxcRom[415] <= 10'b0000100011;
    pxcRom[416] <= 10'b0000001100;
    pxcRom[417] <= 10'b0000000000;
    pxcRom[418] <= 10'b0000000000;
    pxcRom[419] <= 10'b0000000000;
    pxcRom[420] <= 10'b0000000000;
    pxcRom[421] <= 10'b0000000000;
    pxcRom[422] <= 10'b0000000000;
    pxcRom[423] <= 10'b0000000000;
    pxcRom[424] <= 10'b0000000101;
    pxcRom[425] <= 10'b0000011100;
    pxcRom[426] <= 10'b0000111001;
    pxcRom[427] <= 10'b0001011100;
    pxcRom[428] <= 10'b0001100100;
    pxcRom[429] <= 10'b0001000100;
    pxcRom[430] <= 10'b0000100101;
    pxcRom[431] <= 10'b0000001111;
    pxcRom[432] <= 10'b0000000101;
    pxcRom[433] <= 10'b0000000010;
    pxcRom[434] <= 10'b0000000001;
    pxcRom[435] <= 10'b0000000010;
    pxcRom[436] <= 10'b0000000101;
    pxcRom[437] <= 10'b0000001101;
    pxcRom[438] <= 10'b0000011101;
    pxcRom[439] <= 10'b0000110101;
    pxcRom[440] <= 10'b0001010001;
    pxcRom[441] <= 10'b0001010001;
    pxcRom[442] <= 10'b0000111010;
    pxcRom[443] <= 10'b0000011110;
    pxcRom[444] <= 10'b0000001010;
    pxcRom[445] <= 10'b0000000000;
    pxcRom[446] <= 10'b0000000000;
    pxcRom[447] <= 10'b0000000000;
    pxcRom[448] <= 10'b0000000000;
    pxcRom[449] <= 10'b0000000000;
    pxcRom[450] <= 10'b0000000000;
    pxcRom[451] <= 10'b0000000000;
    pxcRom[452] <= 10'b0000000111;
    pxcRom[453] <= 10'b0000100010;
    pxcRom[454] <= 10'b0001000001;
    pxcRom[455] <= 10'b0001100011;
    pxcRom[456] <= 10'b0001011110;
    pxcRom[457] <= 10'b0000111010;
    pxcRom[458] <= 10'b0000011100;
    pxcRom[459] <= 10'b0000001010;
    pxcRom[460] <= 10'b0000000011;
    pxcRom[461] <= 10'b0000000001;
    pxcRom[462] <= 10'b0000000001;
    pxcRom[463] <= 10'b0000000100;
    pxcRom[464] <= 10'b0000001001;
    pxcRom[465] <= 10'b0000010101;
    pxcRom[466] <= 10'b0000101001;
    pxcRom[467] <= 10'b0001000010;
    pxcRom[468] <= 10'b0001010110;
    pxcRom[469] <= 10'b0001001010;
    pxcRom[470] <= 10'b0000110000;
    pxcRom[471] <= 10'b0000011001;
    pxcRom[472] <= 10'b0000001000;
    pxcRom[473] <= 10'b0000000000;
    pxcRom[474] <= 10'b0000000000;
    pxcRom[475] <= 10'b0000000000;
    pxcRom[476] <= 10'b0000000000;
    pxcRom[477] <= 10'b0000000000;
    pxcRom[478] <= 10'b0000000000;
    pxcRom[479] <= 10'b0000000000;
    pxcRom[480] <= 10'b0000001001;
    pxcRom[481] <= 10'b0000100101;
    pxcRom[482] <= 10'b0001000101;
    pxcRom[483] <= 10'b0001100110;
    pxcRom[484] <= 10'b0001011010;
    pxcRom[485] <= 10'b0000110100;
    pxcRom[486] <= 10'b0000011000;
    pxcRom[487] <= 10'b0000001001;
    pxcRom[488] <= 10'b0000000100;
    pxcRom[489] <= 10'b0000000011;
    pxcRom[490] <= 10'b0000000101;
    pxcRom[491] <= 10'b0000001010;
    pxcRom[492] <= 10'b0000010100;
    pxcRom[493] <= 10'b0000100101;
    pxcRom[494] <= 10'b0000111010;
    pxcRom[495] <= 10'b0001010010;
    pxcRom[496] <= 10'b0001010100;
    pxcRom[497] <= 10'b0000111101;
    pxcRom[498] <= 10'b0000100011;
    pxcRom[499] <= 10'b0000010001;
    pxcRom[500] <= 10'b0000000101;
    pxcRom[501] <= 10'b0000000000;
    pxcRom[502] <= 10'b0000000000;
    pxcRom[503] <= 10'b0000000000;
    pxcRom[504] <= 10'b0000000000;
    pxcRom[505] <= 10'b0000000000;
    pxcRom[506] <= 10'b0000000000;
    pxcRom[507] <= 10'b0000000000;
    pxcRom[508] <= 10'b0000001010;
    pxcRom[509] <= 10'b0000100101;
    pxcRom[510] <= 10'b0001000100;
    pxcRom[511] <= 10'b0001100101;
    pxcRom[512] <= 10'b0001011100;
    pxcRom[513] <= 10'b0000111000;
    pxcRom[514] <= 10'b0000011101;
    pxcRom[515] <= 10'b0000001110;
    pxcRom[516] <= 10'b0000001001;
    pxcRom[517] <= 10'b0000001010;
    pxcRom[518] <= 10'b0000001111;
    pxcRom[519] <= 10'b0000011000;
    pxcRom[520] <= 10'b0000100111;
    pxcRom[521] <= 10'b0000111010;
    pxcRom[522] <= 10'b0001010001;
    pxcRom[523] <= 10'b0001011001;
    pxcRom[524] <= 10'b0001000111;
    pxcRom[525] <= 10'b0000101101;
    pxcRom[526] <= 10'b0000011001;
    pxcRom[527] <= 10'b0000001011;
    pxcRom[528] <= 10'b0000000011;
    pxcRom[529] <= 10'b0000000000;
    pxcRom[530] <= 10'b0000000000;
    pxcRom[531] <= 10'b0000000000;
    pxcRom[532] <= 10'b0000000000;
    pxcRom[533] <= 10'b0000000000;
    pxcRom[534] <= 10'b0000000000;
    pxcRom[535] <= 10'b0000000000;
    pxcRom[536] <= 10'b0000001001;
    pxcRom[537] <= 10'b0000100001;
    pxcRom[538] <= 10'b0000111111;
    pxcRom[539] <= 10'b0001100001;
    pxcRom[540] <= 10'b0001100101;
    pxcRom[541] <= 10'b0001001001;
    pxcRom[542] <= 10'b0000101110;
    pxcRom[543] <= 10'b0000011110;
    pxcRom[544] <= 10'b0000011001;
    pxcRom[545] <= 10'b0000011011;
    pxcRom[546] <= 10'b0000100011;
    pxcRom[547] <= 10'b0000110000;
    pxcRom[548] <= 10'b0001000011;
    pxcRom[549] <= 10'b0001010101;
    pxcRom[550] <= 10'b0001011110;
    pxcRom[551] <= 10'b0001001111;
    pxcRom[552] <= 10'b0000110011;
    pxcRom[553] <= 10'b0000011110;
    pxcRom[554] <= 10'b0000001111;
    pxcRom[555] <= 10'b0000000101;
    pxcRom[556] <= 10'b0000000001;
    pxcRom[557] <= 10'b0000000000;
    pxcRom[558] <= 10'b0000000000;
    pxcRom[559] <= 10'b0000000000;
    pxcRom[560] <= 10'b0000000000;
    pxcRom[561] <= 10'b0000000000;
    pxcRom[562] <= 10'b0000000000;
    pxcRom[563] <= 10'b0000000000;
    pxcRom[564] <= 10'b0000000111;
    pxcRom[565] <= 10'b0000011010;
    pxcRom[566] <= 10'b0000110101;
    pxcRom[567] <= 10'b0001010111;
    pxcRom[568] <= 10'b0001110001;
    pxcRom[569] <= 10'b0001101011;
    pxcRom[570] <= 10'b0001010011;
    pxcRom[571] <= 10'b0001000010;
    pxcRom[572] <= 10'b0000111100;
    pxcRom[573] <= 10'b0000111101;
    pxcRom[574] <= 10'b0001000110;
    pxcRom[575] <= 10'b0001010100;
    pxcRom[576] <= 10'b0001100010;
    pxcRom[577] <= 10'b0001100011;
    pxcRom[578] <= 10'b0001010001;
    pxcRom[579] <= 10'b0000110100;
    pxcRom[580] <= 10'b0000100000;
    pxcRom[581] <= 10'b0000010010;
    pxcRom[582] <= 10'b0000000111;
    pxcRom[583] <= 10'b0000000010;
    pxcRom[584] <= 10'b0000000000;
    pxcRom[585] <= 10'b0000000000;
    pxcRom[586] <= 10'b0000000000;
    pxcRom[587] <= 10'b0000000000;
    pxcRom[588] <= 10'b0000000000;
    pxcRom[589] <= 10'b0000000000;
    pxcRom[590] <= 10'b0000000000;
    pxcRom[591] <= 10'b0000000000;
    pxcRom[592] <= 10'b0000000101;
    pxcRom[593] <= 10'b0000010001;
    pxcRom[594] <= 10'b0000100110;
    pxcRom[595] <= 10'b0001000011;
    pxcRom[596] <= 10'b0001101000;
    pxcRom[597] <= 10'b0010001000;
    pxcRom[598] <= 10'b0010001011;
    pxcRom[599] <= 10'b0001111101;
    pxcRom[600] <= 10'b0001110011;
    pxcRom[601] <= 10'b0001110000;
    pxcRom[602] <= 10'b0001110011;
    pxcRom[603] <= 10'b0001110100;
    pxcRom[604] <= 10'b0001100110;
    pxcRom[605] <= 10'b0001001100;
    pxcRom[606] <= 10'b0000110010;
    pxcRom[607] <= 10'b0000011111;
    pxcRom[608] <= 10'b0000010001;
    pxcRom[609] <= 10'b0000001000;
    pxcRom[610] <= 10'b0000000011;
    pxcRom[611] <= 10'b0000000000;
    pxcRom[612] <= 10'b0000000000;
    pxcRom[613] <= 10'b0000000000;
    pxcRom[614] <= 10'b0000000000;
    pxcRom[615] <= 10'b0000000000;
    pxcRom[616] <= 10'b0000000000;
    pxcRom[617] <= 10'b0000000000;
    pxcRom[618] <= 10'b0000000000;
    pxcRom[619] <= 10'b0000000000;
    pxcRom[620] <= 10'b0000000010;
    pxcRom[621] <= 10'b0000001001;
    pxcRom[622] <= 10'b0000010101;
    pxcRom[623] <= 10'b0000101001;
    pxcRom[624] <= 10'b0001000100;
    pxcRom[625] <= 10'b0001100101;
    pxcRom[626] <= 10'b0010000100;
    pxcRom[627] <= 10'b0010001111;
    pxcRom[628] <= 10'b0010001100;
    pxcRom[629] <= 10'b0010000010;
    pxcRom[630] <= 10'b0001110010;
    pxcRom[631] <= 10'b0001011001;
    pxcRom[632] <= 10'b0001000000;
    pxcRom[633] <= 10'b0000101010;
    pxcRom[634] <= 10'b0000011001;
    pxcRom[635] <= 10'b0000001110;
    pxcRom[636] <= 10'b0000000110;
    pxcRom[637] <= 10'b0000000010;
    pxcRom[638] <= 10'b0000000000;
    pxcRom[639] <= 10'b0000000000;
    pxcRom[640] <= 10'b0000000000;
    pxcRom[641] <= 10'b0000000000;
    pxcRom[642] <= 10'b0000000000;
    pxcRom[643] <= 10'b0000000000;
    pxcRom[644] <= 10'b0000000000;
    pxcRom[645] <= 10'b0000000000;
    pxcRom[646] <= 10'b0000000000;
    pxcRom[647] <= 10'b0000000000;
    pxcRom[648] <= 10'b0000000000;
    pxcRom[649] <= 10'b0000000010;
    pxcRom[650] <= 10'b0000001000;
    pxcRom[651] <= 10'b0000010010;
    pxcRom[652] <= 10'b0000100000;
    pxcRom[653] <= 10'b0000110010;
    pxcRom[654] <= 10'b0001000100;
    pxcRom[655] <= 10'b0001010000;
    pxcRom[656] <= 10'b0001010010;
    pxcRom[657] <= 10'b0001001010;
    pxcRom[658] <= 10'b0000111001;
    pxcRom[659] <= 10'b0000101001;
    pxcRom[660] <= 10'b0000011100;
    pxcRom[661] <= 10'b0000010001;
    pxcRom[662] <= 10'b0000001001;
    pxcRom[663] <= 10'b0000000100;
    pxcRom[664] <= 10'b0000000001;
    pxcRom[665] <= 10'b0000000000;
    pxcRom[666] <= 10'b0000000000;
    pxcRom[667] <= 10'b0000000000;
    pxcRom[668] <= 10'b0000000000;
    pxcRom[669] <= 10'b0000000000;
    pxcRom[670] <= 10'b0000000000;
    pxcRom[671] <= 10'b0000000000;
    pxcRom[672] <= 10'b0000000000;
    pxcRom[673] <= 10'b0000000000;
    pxcRom[674] <= 10'b0000000000;
    pxcRom[675] <= 10'b0000000000;
    pxcRom[676] <= 10'b0000000000;
    pxcRom[677] <= 10'b0000000000;
    pxcRom[678] <= 10'b0000000001;
    pxcRom[679] <= 10'b0000000010;
    pxcRom[680] <= 10'b0000000101;
    pxcRom[681] <= 10'b0000001000;
    pxcRom[682] <= 10'b0000001011;
    pxcRom[683] <= 10'b0000001101;
    pxcRom[684] <= 10'b0000001110;
    pxcRom[685] <= 10'b0000001101;
    pxcRom[686] <= 10'b0000001011;
    pxcRom[687] <= 10'b0000001000;
    pxcRom[688] <= 10'b0000000101;
    pxcRom[689] <= 10'b0000000011;
    pxcRom[690] <= 10'b0000000001;
    pxcRom[691] <= 10'b0000000000;
    pxcRom[692] <= 10'b0000000000;
    pxcRom[693] <= 10'b0000000000;
    pxcRom[694] <= 10'b0000000000;
    pxcRom[695] <= 10'b0000000000;
    pxcRom[696] <= 10'b0000000000;
    pxcRom[697] <= 10'b0000000000;
    pxcRom[698] <= 10'b0000000000;
    pxcRom[699] <= 10'b0000000000;
    pxcRom[700] <= 10'b0000000000;
    pxcRom[701] <= 10'b0000000000;
    pxcRom[702] <= 10'b0000000000;
    pxcRom[703] <= 10'b0000000000;
    pxcRom[704] <= 10'b0000000000;
    pxcRom[705] <= 10'b0000000000;
    pxcRom[706] <= 10'b0000000000;
    pxcRom[707] <= 10'b0000000000;
    pxcRom[708] <= 10'b0000000000;
    pxcRom[709] <= 10'b0000000000;
    pxcRom[710] <= 10'b0000000000;
    pxcRom[711] <= 10'b0000000000;
    pxcRom[712] <= 10'b0000000000;
    pxcRom[713] <= 10'b0000000000;
    pxcRom[714] <= 10'b0000000000;
    pxcRom[715] <= 10'b0000000000;
    pxcRom[716] <= 10'b0000000000;
    pxcRom[717] <= 10'b0000000000;
    pxcRom[718] <= 10'b0000000000;
    pxcRom[719] <= 10'b0000000000;
    pxcRom[720] <= 10'b0000000000;
    pxcRom[721] <= 10'b0000000000;
    pxcRom[722] <= 10'b0000000000;
    pxcRom[723] <= 10'b0000000000;
    pxcRom[724] <= 10'b0000000000;
    pxcRom[725] <= 10'b0000000000;
    pxcRom[726] <= 10'b0000000000;
    pxcRom[727] <= 10'b0000000000;
    pxcRom[728] <= 10'b0000000000;
    pxcRom[729] <= 10'b0000000000;
    pxcRom[730] <= 10'b0000000000;
    pxcRom[731] <= 10'b0000000000;
    pxcRom[732] <= 10'b0000000000;
    pxcRom[733] <= 10'b0000000000;
    pxcRom[734] <= 10'b0000000000;
    pxcRom[735] <= 10'b0000000000;
    pxcRom[736] <= 10'b0000000000;
    pxcRom[737] <= 10'b0000000000;
    pxcRom[738] <= 10'b0000000000;
    pxcRom[739] <= 10'b0000000000;
    pxcRom[740] <= 10'b0000000000;
    pxcRom[741] <= 10'b0000000000;
    pxcRom[742] <= 10'b0000000000;
    pxcRom[743] <= 10'b0000000000;
    pxcRom[744] <= 10'b0000000000;
    pxcRom[745] <= 10'b0000000000;
    pxcRom[746] <= 10'b0000000000;
    pxcRom[747] <= 10'b0000000000;
    pxcRom[748] <= 10'b0000000000;
    pxcRom[749] <= 10'b0000000000;
    pxcRom[750] <= 10'b0000000000;
    pxcRom[751] <= 10'b0000000000;
    pxcRom[752] <= 10'b0000000000;
    pxcRom[753] <= 10'b0000000000;
    pxcRom[754] <= 10'b0000000000;
    pxcRom[755] <= 10'b0000000000;
    pxcRom[756] <= 10'b0000000000;
    pxcRom[757] <= 10'b0000000000;
    pxcRom[758] <= 10'b0000000000;
    pxcRom[759] <= 10'b0000000000;
    pxcRom[760] <= 10'b0000000000;
    pxcRom[761] <= 10'b0000000000;
    pxcRom[762] <= 10'b0000000000;
    pxcRom[763] <= 10'b0000000000;
    pxcRom[764] <= 10'b0000000000;
    pxcRom[765] <= 10'b0000000000;
    pxcRom[766] <= 10'b0000000000;
    pxcRom[767] <= 10'b0000000000;
    pxcRom[768] <= 10'b0000000000;
    pxcRom[769] <= 10'b0000000000;
    pxcRom[770] <= 10'b0000000000;
    pxcRom[771] <= 10'b0000000000;
    pxcRom[772] <= 10'b0000000000;
    pxcRom[773] <= 10'b0000000000;
    pxcRom[774] <= 10'b0000000000;
    pxcRom[775] <= 10'b0000000000;
    pxcRom[776] <= 10'b0000000000;
    pxcRom[777] <= 10'b0000000000;
    pxcRom[778] <= 10'b0000000000;
    pxcRom[779] <= 10'b0000000000;
    pxcRom[780] <= 10'b0000000000;
    pxcRom[781] <= 10'b0000000000;
    pxcRom[782] <= 10'b0000000000;
    pxcRom[783] <= 10'b0000000000;
    pxcRom[784] <= 10'b0000000000;
    pxcRom[785] <= 10'b0000000000;
    pxcRom[786] <= 10'b0000000000;
    pxcRom[787] <= 10'b0000000000;
    pxcRom[788] <= 10'b0000000000;
    pxcRom[789] <= 10'b0000000000;
    pxcRom[790] <= 10'b0000000000;
    pxcRom[791] <= 10'b0000000000;
    pxcRom[792] <= 10'b0000000000;
    pxcRom[793] <= 10'b0000000000;
    pxcRom[794] <= 10'b0000000000;
    pxcRom[795] <= 10'b0000000000;
    pxcRom[796] <= 10'b0000000000;
    pxcRom[797] <= 10'b0000000000;
    pxcRom[798] <= 10'b0000000000;
    pxcRom[799] <= 10'b0000000000;
    pxcRom[800] <= 10'b0000000000;
    pxcRom[801] <= 10'b0000000000;
    pxcRom[802] <= 10'b0000000000;
    pxcRom[803] <= 10'b0000000000;
    pxcRom[804] <= 10'b0000000000;
    pxcRom[805] <= 10'b0000000000;
    pxcRom[806] <= 10'b0000000000;
    pxcRom[807] <= 10'b0000000000;
    pxcRom[808] <= 10'b0000000000;
    pxcRom[809] <= 10'b0000000000;
    pxcRom[810] <= 10'b0000000000;
    pxcRom[811] <= 10'b0000000000;
    pxcRom[812] <= 10'b0000000000;
    pxcRom[813] <= 10'b0000000000;
    pxcRom[814] <= 10'b0000000000;
    pxcRom[815] <= 10'b0000000000;
    pxcRom[816] <= 10'b0000000000;
    pxcRom[817] <= 10'b0000000000;
    pxcRom[818] <= 10'b0000000000;
    pxcRom[819] <= 10'b0000000000;
    pxcRom[820] <= 10'b0000000000;
    pxcRom[821] <= 10'b0000000000;
    pxcRom[822] <= 10'b0000000000;
    pxcRom[823] <= 10'b0000000000;
    pxcRom[824] <= 10'b0000000000;
    pxcRom[825] <= 10'b0000000000;
    pxcRom[826] <= 10'b0000000000;
    pxcRom[827] <= 10'b0000000000;
    pxcRom[828] <= 10'b0000000000;
    pxcRom[829] <= 10'b0000000000;
    pxcRom[830] <= 10'b0000000000;
    pxcRom[831] <= 10'b0000000000;
    pxcRom[832] <= 10'b0000000000;
    pxcRom[833] <= 10'b0000000000;
    pxcRom[834] <= 10'b0000000000;
    pxcRom[835] <= 10'b0000000000;
    pxcRom[836] <= 10'b0000000000;
    pxcRom[837] <= 10'b0000000000;
    pxcRom[838] <= 10'b0000000000;
    pxcRom[839] <= 10'b0000000000;
    pxcRom[840] <= 10'b0000000000;
    pxcRom[841] <= 10'b0000000000;
    pxcRom[842] <= 10'b0000000000;
    pxcRom[843] <= 10'b0000000000;
    pxcRom[844] <= 10'b0000000000;
    pxcRom[845] <= 10'b0000000000;
    pxcRom[846] <= 10'b0000000000;
    pxcRom[847] <= 10'b0000000000;
    pxcRom[848] <= 10'b0000000000;
    pxcRom[849] <= 10'b0000000000;
    pxcRom[850] <= 10'b0000000000;
    pxcRom[851] <= 10'b0000000000;
    pxcRom[852] <= 10'b0000000000;
    pxcRom[853] <= 10'b0000000000;
    pxcRom[854] <= 10'b0000000000;
    pxcRom[855] <= 10'b0000000000;
    pxcRom[856] <= 10'b0000000000;
    pxcRom[857] <= 10'b0000000000;
    pxcRom[858] <= 10'b0000000000;
    pxcRom[859] <= 10'b0000000000;
    pxcRom[860] <= 10'b0000000000;
    pxcRom[861] <= 10'b0000000000;
    pxcRom[862] <= 10'b0000000000;
    pxcRom[863] <= 10'b0000000000;
    pxcRom[864] <= 10'b0000000000;
    pxcRom[865] <= 10'b0000000000;
    pxcRom[866] <= 10'b0000000000;
    pxcRom[867] <= 10'b0000000000;
    pxcRom[868] <= 10'b0000000000;
    pxcRom[869] <= 10'b0000000000;
    pxcRom[870] <= 10'b0000000000;
    pxcRom[871] <= 10'b0000000000;
    pxcRom[872] <= 10'b0000000000;
    pxcRom[873] <= 10'b0000000000;
    pxcRom[874] <= 10'b0000000000;
    pxcRom[875] <= 10'b0000000000;
    pxcRom[876] <= 10'b0000000000;
    pxcRom[877] <= 10'b0000000000;
    pxcRom[878] <= 10'b0000000000;
    pxcRom[879] <= 10'b0000000000;
    pxcRom[880] <= 10'b0000000000;
    pxcRom[881] <= 10'b0000000000;
    pxcRom[882] <= 10'b0000000000;
    pxcRom[883] <= 10'b0000000000;
    pxcRom[884] <= 10'b0000000000;
    pxcRom[885] <= 10'b0000000000;
    pxcRom[886] <= 10'b0000000000;
    pxcRom[887] <= 10'b0000000000;
    pxcRom[888] <= 10'b0000000000;
    pxcRom[889] <= 10'b0000000000;
    pxcRom[890] <= 10'b0000000000;
    pxcRom[891] <= 10'b0000000000;
    pxcRom[892] <= 10'b0000000000;
    pxcRom[893] <= 10'b0000000000;
    pxcRom[894] <= 10'b0000000000;
    pxcRom[895] <= 10'b0000000000;
    pxcRom[896] <= 10'b0000000000;
    pxcRom[897] <= 10'b0000000000;
    pxcRom[898] <= 10'b0000000000;
    pxcRom[899] <= 10'b0000000000;
    pxcRom[900] <= 10'b0000000000;
    pxcRom[901] <= 10'b0000000000;
    pxcRom[902] <= 10'b0000000000;
    pxcRom[903] <= 10'b0000000000;
    pxcRom[904] <= 10'b0000000000;
    pxcRom[905] <= 10'b0000000000;
    pxcRom[906] <= 10'b0000000000;
    pxcRom[907] <= 10'b0000000010;
    pxcRom[908] <= 10'b0000000110;
    pxcRom[909] <= 10'b0000001011;
    pxcRom[910] <= 10'b0000010000;
    pxcRom[911] <= 10'b0000010011;
    pxcRom[912] <= 10'b0000010010;
    pxcRom[913] <= 10'b0000010001;
    pxcRom[914] <= 10'b0000001110;
    pxcRom[915] <= 10'b0000001011;
    pxcRom[916] <= 10'b0000000111;
    pxcRom[917] <= 10'b0000000011;
    pxcRom[918] <= 10'b0000000001;
    pxcRom[919] <= 10'b0000000000;
    pxcRom[920] <= 10'b0000000000;
    pxcRom[921] <= 10'b0000000000;
    pxcRom[922] <= 10'b0000000000;
    pxcRom[923] <= 10'b0000000000;
    pxcRom[924] <= 10'b0000000000;
    pxcRom[925] <= 10'b0000000000;
    pxcRom[926] <= 10'b0000000000;
    pxcRom[927] <= 10'b0000000000;
    pxcRom[928] <= 10'b0000000000;
    pxcRom[929] <= 10'b0000000000;
    pxcRom[930] <= 10'b0000000000;
    pxcRom[931] <= 10'b0000000000;
    pxcRom[932] <= 10'b0000000000;
    pxcRom[933] <= 10'b0000000000;
    pxcRom[934] <= 10'b0000000001;
    pxcRom[935] <= 10'b0000000100;
    pxcRom[936] <= 10'b0000001010;
    pxcRom[937] <= 10'b0000010101;
    pxcRom[938] <= 10'b0000100000;
    pxcRom[939] <= 10'b0000101000;
    pxcRom[940] <= 10'b0000101001;
    pxcRom[941] <= 10'b0000100100;
    pxcRom[942] <= 10'b0000011100;
    pxcRom[943] <= 10'b0000010100;
    pxcRom[944] <= 10'b0000001100;
    pxcRom[945] <= 10'b0000000110;
    pxcRom[946] <= 10'b0000000010;
    pxcRom[947] <= 10'b0000000001;
    pxcRom[948] <= 10'b0000000000;
    pxcRom[949] <= 10'b0000000000;
    pxcRom[950] <= 10'b0000000000;
    pxcRom[951] <= 10'b0000000000;
    pxcRom[952] <= 10'b0000000000;
    pxcRom[953] <= 10'b0000000000;
    pxcRom[954] <= 10'b0000000000;
    pxcRom[955] <= 10'b0000000000;
    pxcRom[956] <= 10'b0000000000;
    pxcRom[957] <= 10'b0000000000;
    pxcRom[958] <= 10'b0000000000;
    pxcRom[959] <= 10'b0000000000;
    pxcRom[960] <= 10'b0000000000;
    pxcRom[961] <= 10'b0000000000;
    pxcRom[962] <= 10'b0000000001;
    pxcRom[963] <= 10'b0000000100;
    pxcRom[964] <= 10'b0000001011;
    pxcRom[965] <= 10'b0000011000;
    pxcRom[966] <= 10'b0000101000;
    pxcRom[967] <= 10'b0000110100;
    pxcRom[968] <= 10'b0000110110;
    pxcRom[969] <= 10'b0000101101;
    pxcRom[970] <= 10'b0000100001;
    pxcRom[971] <= 10'b0000010101;
    pxcRom[972] <= 10'b0000001100;
    pxcRom[973] <= 10'b0000000110;
    pxcRom[974] <= 10'b0000000010;
    pxcRom[975] <= 10'b0000000000;
    pxcRom[976] <= 10'b0000000000;
    pxcRom[977] <= 10'b0000000000;
    pxcRom[978] <= 10'b0000000000;
    pxcRom[979] <= 10'b0000000000;
    pxcRom[980] <= 10'b0000000000;
    pxcRom[981] <= 10'b0000000000;
    pxcRom[982] <= 10'b0000000000;
    pxcRom[983] <= 10'b0000000000;
    pxcRom[984] <= 10'b0000000000;
    pxcRom[985] <= 10'b0000000000;
    pxcRom[986] <= 10'b0000000000;
    pxcRom[987] <= 10'b0000000000;
    pxcRom[988] <= 10'b0000000000;
    pxcRom[989] <= 10'b0000000000;
    pxcRom[990] <= 10'b0000000001;
    pxcRom[991] <= 10'b0000000100;
    pxcRom[992] <= 10'b0000001100;
    pxcRom[993] <= 10'b0000011011;
    pxcRom[994] <= 10'b0000101111;
    pxcRom[995] <= 10'b0001000010;
    pxcRom[996] <= 10'b0001000000;
    pxcRom[997] <= 10'b0000110001;
    pxcRom[998] <= 10'b0000100000;
    pxcRom[999] <= 10'b0000010011;
    pxcRom[1000] <= 10'b0000001010;
    pxcRom[1001] <= 10'b0000000100;
    pxcRom[1002] <= 10'b0000000001;
    pxcRom[1003] <= 10'b0000000000;
    pxcRom[1004] <= 10'b0000000000;
    pxcRom[1005] <= 10'b0000000000;
    pxcRom[1006] <= 10'b0000000000;
    pxcRom[1007] <= 10'b0000000000;
    pxcRom[1008] <= 10'b0000000000;
    pxcRom[1009] <= 10'b0000000000;
    pxcRom[1010] <= 10'b0000000000;
    pxcRom[1011] <= 10'b0000000000;
    pxcRom[1012] <= 10'b0000000000;
    pxcRom[1013] <= 10'b0000000000;
    pxcRom[1014] <= 10'b0000000000;
    pxcRom[1015] <= 10'b0000000000;
    pxcRom[1016] <= 10'b0000000000;
    pxcRom[1017] <= 10'b0000000000;
    pxcRom[1018] <= 10'b0000000001;
    pxcRom[1019] <= 10'b0000000100;
    pxcRom[1020] <= 10'b0000001100;
    pxcRom[1021] <= 10'b0000011101;
    pxcRom[1022] <= 10'b0000111000;
    pxcRom[1023] <= 10'b0001010010;
    pxcRom[1024] <= 10'b0001001100;
    pxcRom[1025] <= 10'b0000110010;
    pxcRom[1026] <= 10'b0000011100;
    pxcRom[1027] <= 10'b0000001111;
    pxcRom[1028] <= 10'b0000000110;
    pxcRom[1029] <= 10'b0000000010;
    pxcRom[1030] <= 10'b0000000000;
    pxcRom[1031] <= 10'b0000000000;
    pxcRom[1032] <= 10'b0000000000;
    pxcRom[1033] <= 10'b0000000000;
    pxcRom[1034] <= 10'b0000000000;
    pxcRom[1035] <= 10'b0000000000;
    pxcRom[1036] <= 10'b0000000000;
    pxcRom[1037] <= 10'b0000000000;
    pxcRom[1038] <= 10'b0000000000;
    pxcRom[1039] <= 10'b0000000000;
    pxcRom[1040] <= 10'b0000000000;
    pxcRom[1041] <= 10'b0000000000;
    pxcRom[1042] <= 10'b0000000000;
    pxcRom[1043] <= 10'b0000000000;
    pxcRom[1044] <= 10'b0000000000;
    pxcRom[1045] <= 10'b0000000000;
    pxcRom[1046] <= 10'b0000000001;
    pxcRom[1047] <= 10'b0000000011;
    pxcRom[1048] <= 10'b0000001100;
    pxcRom[1049] <= 10'b0000100001;
    pxcRom[1050] <= 10'b0001001000;
    pxcRom[1051] <= 10'b0001101111;
    pxcRom[1052] <= 10'b0001010100;
    pxcRom[1053] <= 10'b0000101110;
    pxcRom[1054] <= 10'b0000011000;
    pxcRom[1055] <= 10'b0000001010;
    pxcRom[1056] <= 10'b0000000011;
    pxcRom[1057] <= 10'b0000000001;
    pxcRom[1058] <= 10'b0000000000;
    pxcRom[1059] <= 10'b0000000000;
    pxcRom[1060] <= 10'b0000000000;
    pxcRom[1061] <= 10'b0000000000;
    pxcRom[1062] <= 10'b0000000000;
    pxcRom[1063] <= 10'b0000000000;
    pxcRom[1064] <= 10'b0000000000;
    pxcRom[1065] <= 10'b0000000000;
    pxcRom[1066] <= 10'b0000000000;
    pxcRom[1067] <= 10'b0000000000;
    pxcRom[1068] <= 10'b0000000000;
    pxcRom[1069] <= 10'b0000000000;
    pxcRom[1070] <= 10'b0000000000;
    pxcRom[1071] <= 10'b0000000000;
    pxcRom[1072] <= 10'b0000000000;
    pxcRom[1073] <= 10'b0000000000;
    pxcRom[1074] <= 10'b0000000001;
    pxcRom[1075] <= 10'b0000000011;
    pxcRom[1076] <= 10'b0000001100;
    pxcRom[1077] <= 10'b0000100111;
    pxcRom[1078] <= 10'b0001100011;
    pxcRom[1079] <= 10'b0010010111;
    pxcRom[1080] <= 10'b0001010101;
    pxcRom[1081] <= 10'b0000100111;
    pxcRom[1082] <= 10'b0000010001;
    pxcRom[1083] <= 10'b0000000110;
    pxcRom[1084] <= 10'b0000000001;
    pxcRom[1085] <= 10'b0000000000;
    pxcRom[1086] <= 10'b0000000000;
    pxcRom[1087] <= 10'b0000000000;
    pxcRom[1088] <= 10'b0000000000;
    pxcRom[1089] <= 10'b0000000000;
    pxcRom[1090] <= 10'b0000000000;
    pxcRom[1091] <= 10'b0000000000;
    pxcRom[1092] <= 10'b0000000000;
    pxcRom[1093] <= 10'b0000000000;
    pxcRom[1094] <= 10'b0000000000;
    pxcRom[1095] <= 10'b0000000000;
    pxcRom[1096] <= 10'b0000000000;
    pxcRom[1097] <= 10'b0000000000;
    pxcRom[1098] <= 10'b0000000000;
    pxcRom[1099] <= 10'b0000000000;
    pxcRom[1100] <= 10'b0000000000;
    pxcRom[1101] <= 10'b0000000000;
    pxcRom[1102] <= 10'b0000000001;
    pxcRom[1103] <= 10'b0000000010;
    pxcRom[1104] <= 10'b0000001101;
    pxcRom[1105] <= 10'b0000110100;
    pxcRom[1106] <= 10'b0010010101;
    pxcRom[1107] <= 10'b0010111011;
    pxcRom[1108] <= 10'b0001010000;
    pxcRom[1109] <= 10'b0000011111;
    pxcRom[1110] <= 10'b0000001010;
    pxcRom[1111] <= 10'b0000000010;
    pxcRom[1112] <= 10'b0000000000;
    pxcRom[1113] <= 10'b0000000000;
    pxcRom[1114] <= 10'b0000000000;
    pxcRom[1115] <= 10'b0000000000;
    pxcRom[1116] <= 10'b0000000000;
    pxcRom[1117] <= 10'b0000000000;
    pxcRom[1118] <= 10'b0000000000;
    pxcRom[1119] <= 10'b0000000000;
    pxcRom[1120] <= 10'b0000000000;
    pxcRom[1121] <= 10'b0000000000;
    pxcRom[1122] <= 10'b0000000000;
    pxcRom[1123] <= 10'b0000000000;
    pxcRom[1124] <= 10'b0000000000;
    pxcRom[1125] <= 10'b0000000000;
    pxcRom[1126] <= 10'b0000000000;
    pxcRom[1127] <= 10'b0000000000;
    pxcRom[1128] <= 10'b0000000000;
    pxcRom[1129] <= 10'b0000000000;
    pxcRom[1130] <= 10'b0000000001;
    pxcRom[1131] <= 10'b0000000010;
    pxcRom[1132] <= 10'b0000001111;
    pxcRom[1133] <= 10'b0001001111;
    pxcRom[1134] <= 10'b0011101100;
    pxcRom[1135] <= 10'b0011001110;
    pxcRom[1136] <= 10'b0001001001;
    pxcRom[1137] <= 10'b0000010100;
    pxcRom[1138] <= 10'b0000000101;
    pxcRom[1139] <= 10'b0000000000;
    pxcRom[1140] <= 10'b0000000000;
    pxcRom[1141] <= 10'b0000000000;
    pxcRom[1142] <= 10'b0000000000;
    pxcRom[1143] <= 10'b0000000000;
    pxcRom[1144] <= 10'b0000000000;
    pxcRom[1145] <= 10'b0000000000;
    pxcRom[1146] <= 10'b0000000000;
    pxcRom[1147] <= 10'b0000000000;
    pxcRom[1148] <= 10'b0000000000;
    pxcRom[1149] <= 10'b0000000000;
    pxcRom[1150] <= 10'b0000000000;
    pxcRom[1151] <= 10'b0000000000;
    pxcRom[1152] <= 10'b0000000000;
    pxcRom[1153] <= 10'b0000000000;
    pxcRom[1154] <= 10'b0000000000;
    pxcRom[1155] <= 10'b0000000000;
    pxcRom[1156] <= 10'b0000000000;
    pxcRom[1157] <= 10'b0000000000;
    pxcRom[1158] <= 10'b0000000000;
    pxcRom[1159] <= 10'b0000000011;
    pxcRom[1160] <= 10'b0000010110;
    pxcRom[1161] <= 10'b0001111111;
    pxcRom[1162] <= 10'b0100101011;
    pxcRom[1163] <= 10'b0011001101;
    pxcRom[1164] <= 10'b0000111010;
    pxcRom[1165] <= 10'b0000001011;
    pxcRom[1166] <= 10'b0000000001;
    pxcRom[1167] <= 10'b0000000000;
    pxcRom[1168] <= 10'b0000000000;
    pxcRom[1169] <= 10'b0000000000;
    pxcRom[1170] <= 10'b0000000000;
    pxcRom[1171] <= 10'b0000000000;
    pxcRom[1172] <= 10'b0000000000;
    pxcRom[1173] <= 10'b0000000000;
    pxcRom[1174] <= 10'b0000000000;
    pxcRom[1175] <= 10'b0000000000;
    pxcRom[1176] <= 10'b0000000000;
    pxcRom[1177] <= 10'b0000000000;
    pxcRom[1178] <= 10'b0000000000;
    pxcRom[1179] <= 10'b0000000000;
    pxcRom[1180] <= 10'b0000000000;
    pxcRom[1181] <= 10'b0000000000;
    pxcRom[1182] <= 10'b0000000000;
    pxcRom[1183] <= 10'b0000000000;
    pxcRom[1184] <= 10'b0000000000;
    pxcRom[1185] <= 10'b0000000000;
    pxcRom[1186] <= 10'b0000000001;
    pxcRom[1187] <= 10'b0000000101;
    pxcRom[1188] <= 10'b0000100100;
    pxcRom[1189] <= 10'b0010101100;
    pxcRom[1190] <= 10'b0100111001;
    pxcRom[1191] <= 10'b0010110100;
    pxcRom[1192] <= 10'b0000100111;
    pxcRom[1193] <= 10'b0000000101;
    pxcRom[1194] <= 10'b0000000000;
    pxcRom[1195] <= 10'b0000000000;
    pxcRom[1196] <= 10'b0000000000;
    pxcRom[1197] <= 10'b0000000000;
    pxcRom[1198] <= 10'b0000000000;
    pxcRom[1199] <= 10'b0000000000;
    pxcRom[1200] <= 10'b0000000000;
    pxcRom[1201] <= 10'b0000000000;
    pxcRom[1202] <= 10'b0000000000;
    pxcRom[1203] <= 10'b0000000000;
    pxcRom[1204] <= 10'b0000000000;
    pxcRom[1205] <= 10'b0000000000;
    pxcRom[1206] <= 10'b0000000000;
    pxcRom[1207] <= 10'b0000000000;
    pxcRom[1208] <= 10'b0000000000;
    pxcRom[1209] <= 10'b0000000000;
    pxcRom[1210] <= 10'b0000000000;
    pxcRom[1211] <= 10'b0000000000;
    pxcRom[1212] <= 10'b0000000000;
    pxcRom[1213] <= 10'b0000000000;
    pxcRom[1214] <= 10'b0000000010;
    pxcRom[1215] <= 10'b0000001011;
    pxcRom[1216] <= 10'b0000110111;
    pxcRom[1217] <= 10'b0011000101;
    pxcRom[1218] <= 10'b0100101101;
    pxcRom[1219] <= 10'b0010000010;
    pxcRom[1220] <= 10'b0000011000;
    pxcRom[1221] <= 10'b0000000010;
    pxcRom[1222] <= 10'b0000000000;
    pxcRom[1223] <= 10'b0000000000;
    pxcRom[1224] <= 10'b0000000000;
    pxcRom[1225] <= 10'b0000000000;
    pxcRom[1226] <= 10'b0000000000;
    pxcRom[1227] <= 10'b0000000000;
    pxcRom[1228] <= 10'b0000000000;
    pxcRom[1229] <= 10'b0000000000;
    pxcRom[1230] <= 10'b0000000000;
    pxcRom[1231] <= 10'b0000000000;
    pxcRom[1232] <= 10'b0000000000;
    pxcRom[1233] <= 10'b0000000000;
    pxcRom[1234] <= 10'b0000000000;
    pxcRom[1235] <= 10'b0000000000;
    pxcRom[1236] <= 10'b0000000000;
    pxcRom[1237] <= 10'b0000000000;
    pxcRom[1238] <= 10'b0000000000;
    pxcRom[1239] <= 10'b0000000000;
    pxcRom[1240] <= 10'b0000000000;
    pxcRom[1241] <= 10'b0000000001;
    pxcRom[1242] <= 10'b0000000101;
    pxcRom[1243] <= 10'b0000010101;
    pxcRom[1244] <= 10'b0001000100;
    pxcRom[1245] <= 10'b0011000001;
    pxcRom[1246] <= 10'b0011100100;
    pxcRom[1247] <= 10'b0001010010;
    pxcRom[1248] <= 10'b0000010000;
    pxcRom[1249] <= 10'b0000000010;
    pxcRom[1250] <= 10'b0000000000;
    pxcRom[1251] <= 10'b0000000000;
    pxcRom[1252] <= 10'b0000000000;
    pxcRom[1253] <= 10'b0000000000;
    pxcRom[1254] <= 10'b0000000000;
    pxcRom[1255] <= 10'b0000000000;
    pxcRom[1256] <= 10'b0000000000;
    pxcRom[1257] <= 10'b0000000000;
    pxcRom[1258] <= 10'b0000000000;
    pxcRom[1259] <= 10'b0000000000;
    pxcRom[1260] <= 10'b0000000000;
    pxcRom[1261] <= 10'b0000000000;
    pxcRom[1262] <= 10'b0000000000;
    pxcRom[1263] <= 10'b0000000000;
    pxcRom[1264] <= 10'b0000000000;
    pxcRom[1265] <= 10'b0000000000;
    pxcRom[1266] <= 10'b0000000000;
    pxcRom[1267] <= 10'b0000000000;
    pxcRom[1268] <= 10'b0000000000;
    pxcRom[1269] <= 10'b0000000011;
    pxcRom[1270] <= 10'b0000001011;
    pxcRom[1271] <= 10'b0000100000;
    pxcRom[1272] <= 10'b0001001100;
    pxcRom[1273] <= 10'b0010101111;
    pxcRom[1274] <= 10'b0010010101;
    pxcRom[1275] <= 10'b0000110110;
    pxcRom[1276] <= 10'b0000001101;
    pxcRom[1277] <= 10'b0000000010;
    pxcRom[1278] <= 10'b0000000000;
    pxcRom[1279] <= 10'b0000000000;
    pxcRom[1280] <= 10'b0000000000;
    pxcRom[1281] <= 10'b0000000000;
    pxcRom[1282] <= 10'b0000000000;
    pxcRom[1283] <= 10'b0000000000;
    pxcRom[1284] <= 10'b0000000000;
    pxcRom[1285] <= 10'b0000000000;
    pxcRom[1286] <= 10'b0000000000;
    pxcRom[1287] <= 10'b0000000000;
    pxcRom[1288] <= 10'b0000000000;
    pxcRom[1289] <= 10'b0000000000;
    pxcRom[1290] <= 10'b0000000000;
    pxcRom[1291] <= 10'b0000000000;
    pxcRom[1292] <= 10'b0000000000;
    pxcRom[1293] <= 10'b0000000000;
    pxcRom[1294] <= 10'b0000000000;
    pxcRom[1295] <= 10'b0000000000;
    pxcRom[1296] <= 10'b0000000010;
    pxcRom[1297] <= 10'b0000000111;
    pxcRom[1298] <= 10'b0000010010;
    pxcRom[1299] <= 10'b0000100111;
    pxcRom[1300] <= 10'b0001010000;
    pxcRom[1301] <= 10'b0010001101;
    pxcRom[1302] <= 10'b0001100001;
    pxcRom[1303] <= 10'b0000101001;
    pxcRom[1304] <= 10'b0000001101;
    pxcRom[1305] <= 10'b0000000011;
    pxcRom[1306] <= 10'b0000000000;
    pxcRom[1307] <= 10'b0000000000;
    pxcRom[1308] <= 10'b0000000000;
    pxcRom[1309] <= 10'b0000000000;
    pxcRom[1310] <= 10'b0000000000;
    pxcRom[1311] <= 10'b0000000000;
    pxcRom[1312] <= 10'b0000000000;
    pxcRom[1313] <= 10'b0000000000;
    pxcRom[1314] <= 10'b0000000000;
    pxcRom[1315] <= 10'b0000000000;
    pxcRom[1316] <= 10'b0000000000;
    pxcRom[1317] <= 10'b0000000000;
    pxcRom[1318] <= 10'b0000000000;
    pxcRom[1319] <= 10'b0000000000;
    pxcRom[1320] <= 10'b0000000000;
    pxcRom[1321] <= 10'b0000000000;
    pxcRom[1322] <= 10'b0000000000;
    pxcRom[1323] <= 10'b0000000001;
    pxcRom[1324] <= 10'b0000000100;
    pxcRom[1325] <= 10'b0000001100;
    pxcRom[1326] <= 10'b0000011010;
    pxcRom[1327] <= 10'b0000101110;
    pxcRom[1328] <= 10'b0001001110;
    pxcRom[1329] <= 10'b0001101100;
    pxcRom[1330] <= 10'b0001000111;
    pxcRom[1331] <= 10'b0000100011;
    pxcRom[1332] <= 10'b0000001110;
    pxcRom[1333] <= 10'b0000000100;
    pxcRom[1334] <= 10'b0000000001;
    pxcRom[1335] <= 10'b0000000000;
    pxcRom[1336] <= 10'b0000000000;
    pxcRom[1337] <= 10'b0000000000;
    pxcRom[1338] <= 10'b0000000000;
    pxcRom[1339] <= 10'b0000000000;
    pxcRom[1340] <= 10'b0000000000;
    pxcRom[1341] <= 10'b0000000000;
    pxcRom[1342] <= 10'b0000000000;
    pxcRom[1343] <= 10'b0000000000;
    pxcRom[1344] <= 10'b0000000000;
    pxcRom[1345] <= 10'b0000000000;
    pxcRom[1346] <= 10'b0000000000;
    pxcRom[1347] <= 10'b0000000000;
    pxcRom[1348] <= 10'b0000000000;
    pxcRom[1349] <= 10'b0000000000;
    pxcRom[1350] <= 10'b0000000001;
    pxcRom[1351] <= 10'b0000000011;
    pxcRom[1352] <= 10'b0000001000;
    pxcRom[1353] <= 10'b0000010001;
    pxcRom[1354] <= 10'b0000011111;
    pxcRom[1355] <= 10'b0000110001;
    pxcRom[1356] <= 10'b0001000111;
    pxcRom[1357] <= 10'b0001010010;
    pxcRom[1358] <= 10'b0000111001;
    pxcRom[1359] <= 10'b0000100000;
    pxcRom[1360] <= 10'b0000001111;
    pxcRom[1361] <= 10'b0000000101;
    pxcRom[1362] <= 10'b0000000010;
    pxcRom[1363] <= 10'b0000000001;
    pxcRom[1364] <= 10'b0000000000;
    pxcRom[1365] <= 10'b0000000000;
    pxcRom[1366] <= 10'b0000000000;
    pxcRom[1367] <= 10'b0000000000;
    pxcRom[1368] <= 10'b0000000000;
    pxcRom[1369] <= 10'b0000000000;
    pxcRom[1370] <= 10'b0000000000;
    pxcRom[1371] <= 10'b0000000000;
    pxcRom[1372] <= 10'b0000000000;
    pxcRom[1373] <= 10'b0000000000;
    pxcRom[1374] <= 10'b0000000000;
    pxcRom[1375] <= 10'b0000000000;
    pxcRom[1376] <= 10'b0000000000;
    pxcRom[1377] <= 10'b0000000000;
    pxcRom[1378] <= 10'b0000000010;
    pxcRom[1379] <= 10'b0000000101;
    pxcRom[1380] <= 10'b0000001011;
    pxcRom[1381] <= 10'b0000010101;
    pxcRom[1382] <= 10'b0000100011;
    pxcRom[1383] <= 10'b0000110001;
    pxcRom[1384] <= 10'b0000111110;
    pxcRom[1385] <= 10'b0001000000;
    pxcRom[1386] <= 10'b0000110001;
    pxcRom[1387] <= 10'b0000011110;
    pxcRom[1388] <= 10'b0000010000;
    pxcRom[1389] <= 10'b0000000111;
    pxcRom[1390] <= 10'b0000000010;
    pxcRom[1391] <= 10'b0000000001;
    pxcRom[1392] <= 10'b0000000000;
    pxcRom[1393] <= 10'b0000000000;
    pxcRom[1394] <= 10'b0000000000;
    pxcRom[1395] <= 10'b0000000000;
    pxcRom[1396] <= 10'b0000000000;
    pxcRom[1397] <= 10'b0000000000;
    pxcRom[1398] <= 10'b0000000000;
    pxcRom[1399] <= 10'b0000000000;
    pxcRom[1400] <= 10'b0000000000;
    pxcRom[1401] <= 10'b0000000000;
    pxcRom[1402] <= 10'b0000000000;
    pxcRom[1403] <= 10'b0000000000;
    pxcRom[1404] <= 10'b0000000000;
    pxcRom[1405] <= 10'b0000000001;
    pxcRom[1406] <= 10'b0000000010;
    pxcRom[1407] <= 10'b0000000110;
    pxcRom[1408] <= 10'b0000001110;
    pxcRom[1409] <= 10'b0000010111;
    pxcRom[1410] <= 10'b0000100010;
    pxcRom[1411] <= 10'b0000101100;
    pxcRom[1412] <= 10'b0000110011;
    pxcRom[1413] <= 10'b0000110011;
    pxcRom[1414] <= 10'b0000101011;
    pxcRom[1415] <= 10'b0000011101;
    pxcRom[1416] <= 10'b0000010000;
    pxcRom[1417] <= 10'b0000000111;
    pxcRom[1418] <= 10'b0000000010;
    pxcRom[1419] <= 10'b0000000001;
    pxcRom[1420] <= 10'b0000000000;
    pxcRom[1421] <= 10'b0000000000;
    pxcRom[1422] <= 10'b0000000000;
    pxcRom[1423] <= 10'b0000000000;
    pxcRom[1424] <= 10'b0000000000;
    pxcRom[1425] <= 10'b0000000000;
    pxcRom[1426] <= 10'b0000000000;
    pxcRom[1427] <= 10'b0000000000;
    pxcRom[1428] <= 10'b0000000000;
    pxcRom[1429] <= 10'b0000000000;
    pxcRom[1430] <= 10'b0000000000;
    pxcRom[1431] <= 10'b0000000000;
    pxcRom[1432] <= 10'b0000000000;
    pxcRom[1433] <= 10'b0000000001;
    pxcRom[1434] <= 10'b0000000010;
    pxcRom[1435] <= 10'b0000000110;
    pxcRom[1436] <= 10'b0000001100;
    pxcRom[1437] <= 10'b0000010100;
    pxcRom[1438] <= 10'b0000011100;
    pxcRom[1439] <= 10'b0000100001;
    pxcRom[1440] <= 10'b0000100100;
    pxcRom[1441] <= 10'b0000100101;
    pxcRom[1442] <= 10'b0000100001;
    pxcRom[1443] <= 10'b0000010111;
    pxcRom[1444] <= 10'b0000001101;
    pxcRom[1445] <= 10'b0000000101;
    pxcRom[1446] <= 10'b0000000001;
    pxcRom[1447] <= 10'b0000000000;
    pxcRom[1448] <= 10'b0000000000;
    pxcRom[1449] <= 10'b0000000000;
    pxcRom[1450] <= 10'b0000000000;
    pxcRom[1451] <= 10'b0000000000;
    pxcRom[1452] <= 10'b0000000000;
    pxcRom[1453] <= 10'b0000000000;
    pxcRom[1454] <= 10'b0000000000;
    pxcRom[1455] <= 10'b0000000000;
    pxcRom[1456] <= 10'b0000000000;
    pxcRom[1457] <= 10'b0000000000;
    pxcRom[1458] <= 10'b0000000000;
    pxcRom[1459] <= 10'b0000000000;
    pxcRom[1460] <= 10'b0000000000;
    pxcRom[1461] <= 10'b0000000000;
    pxcRom[1462] <= 10'b0000000000;
    pxcRom[1463] <= 10'b0000000001;
    pxcRom[1464] <= 10'b0000000011;
    pxcRom[1465] <= 10'b0000000101;
    pxcRom[1466] <= 10'b0000000110;
    pxcRom[1467] <= 10'b0000001000;
    pxcRom[1468] <= 10'b0000001000;
    pxcRom[1469] <= 10'b0000001001;
    pxcRom[1470] <= 10'b0000001000;
    pxcRom[1471] <= 10'b0000000110;
    pxcRom[1472] <= 10'b0000000011;
    pxcRom[1473] <= 10'b0000000001;
    pxcRom[1474] <= 10'b0000000000;
    pxcRom[1475] <= 10'b0000000000;
    pxcRom[1476] <= 10'b0000000000;
    pxcRom[1477] <= 10'b0000000000;
    pxcRom[1478] <= 10'b0000000000;
    pxcRom[1479] <= 10'b0000000000;
    pxcRom[1480] <= 10'b0000000000;
    pxcRom[1481] <= 10'b0000000000;
    pxcRom[1482] <= 10'b0000000000;
    pxcRom[1483] <= 10'b0000000000;
    pxcRom[1484] <= 10'b0000000000;
    pxcRom[1485] <= 10'b0000000000;
    pxcRom[1486] <= 10'b0000000000;
    pxcRom[1487] <= 10'b0000000000;
    pxcRom[1488] <= 10'b0000000000;
    pxcRom[1489] <= 10'b0000000000;
    pxcRom[1490] <= 10'b0000000000;
    pxcRom[1491] <= 10'b0000000000;
    pxcRom[1492] <= 10'b0000000000;
    pxcRom[1493] <= 10'b0000000000;
    pxcRom[1494] <= 10'b0000000000;
    pxcRom[1495] <= 10'b0000000000;
    pxcRom[1496] <= 10'b0000000000;
    pxcRom[1497] <= 10'b0000000000;
    pxcRom[1498] <= 10'b0000000000;
    pxcRom[1499] <= 10'b0000000000;
    pxcRom[1500] <= 10'b0000000000;
    pxcRom[1501] <= 10'b0000000000;
    pxcRom[1502] <= 10'b0000000000;
    pxcRom[1503] <= 10'b0000000000;
    pxcRom[1504] <= 10'b0000000000;
    pxcRom[1505] <= 10'b0000000000;
    pxcRom[1506] <= 10'b0000000000;
    pxcRom[1507] <= 10'b0000000000;
    pxcRom[1508] <= 10'b0000000000;
    pxcRom[1509] <= 10'b0000000000;
    pxcRom[1510] <= 10'b0000000000;
    pxcRom[1511] <= 10'b0000000000;
    pxcRom[1512] <= 10'b0000000000;
    pxcRom[1513] <= 10'b0000000000;
    pxcRom[1514] <= 10'b0000000000;
    pxcRom[1515] <= 10'b0000000000;
    pxcRom[1516] <= 10'b0000000000;
    pxcRom[1517] <= 10'b0000000000;
    pxcRom[1518] <= 10'b0000000000;
    pxcRom[1519] <= 10'b0000000000;
    pxcRom[1520] <= 10'b0000000000;
    pxcRom[1521] <= 10'b0000000000;
    pxcRom[1522] <= 10'b0000000000;
    pxcRom[1523] <= 10'b0000000000;
    pxcRom[1524] <= 10'b0000000000;
    pxcRom[1525] <= 10'b0000000000;
    pxcRom[1526] <= 10'b0000000000;
    pxcRom[1527] <= 10'b0000000000;
    pxcRom[1528] <= 10'b0000000000;
    pxcRom[1529] <= 10'b0000000000;
    pxcRom[1530] <= 10'b0000000000;
    pxcRom[1531] <= 10'b0000000000;
    pxcRom[1532] <= 10'b0000000000;
    pxcRom[1533] <= 10'b0000000000;
    pxcRom[1534] <= 10'b0000000000;
    pxcRom[1535] <= 10'b0000000000;
    pxcRom[1536] <= 10'b0000000000;
    pxcRom[1537] <= 10'b0000000000;
    pxcRom[1538] <= 10'b0000000000;
    pxcRom[1539] <= 10'b0000000000;
    pxcRom[1540] <= 10'b0000000000;
    pxcRom[1541] <= 10'b0000000000;
    pxcRom[1542] <= 10'b0000000000;
    pxcRom[1543] <= 10'b0000000000;
    pxcRom[1544] <= 10'b0000000000;
    pxcRom[1545] <= 10'b0000000000;
    pxcRom[1546] <= 10'b0000000000;
    pxcRom[1547] <= 10'b0000000000;
    pxcRom[1548] <= 10'b0000000000;
    pxcRom[1549] <= 10'b0000000000;
    pxcRom[1550] <= 10'b0000000000;
    pxcRom[1551] <= 10'b0000000000;
    pxcRom[1552] <= 10'b0000000000;
    pxcRom[1553] <= 10'b0000000000;
    pxcRom[1554] <= 10'b0000000000;
    pxcRom[1555] <= 10'b0000000000;
    pxcRom[1556] <= 10'b0000000000;
    pxcRom[1557] <= 10'b0000000000;
    pxcRom[1558] <= 10'b0000000000;
    pxcRom[1559] <= 10'b0000000000;
    pxcRom[1560] <= 10'b0000000000;
    pxcRom[1561] <= 10'b0000000000;
    pxcRom[1562] <= 10'b0000000000;
    pxcRom[1563] <= 10'b0000000000;
    pxcRom[1564] <= 10'b0000000000;
    pxcRom[1565] <= 10'b0000000000;
    pxcRom[1566] <= 10'b0000000000;
    pxcRom[1567] <= 10'b0000000000;
    pxcRom[1568] <= 10'b0000000000;
    pxcRom[1569] <= 10'b0000000000;
    pxcRom[1570] <= 10'b0000000000;
    pxcRom[1571] <= 10'b0000000000;
    pxcRom[1572] <= 10'b0000000000;
    pxcRom[1573] <= 10'b0000000000;
    pxcRom[1574] <= 10'b0000000000;
    pxcRom[1575] <= 10'b0000000000;
    pxcRom[1576] <= 10'b0000000000;
    pxcRom[1577] <= 10'b0000000000;
    pxcRom[1578] <= 10'b0000000000;
    pxcRom[1579] <= 10'b0000000000;
    pxcRom[1580] <= 10'b0000000000;
    pxcRom[1581] <= 10'b0000000000;
    pxcRom[1582] <= 10'b0000000000;
    pxcRom[1583] <= 10'b0000000000;
    pxcRom[1584] <= 10'b0000000000;
    pxcRom[1585] <= 10'b0000000000;
    pxcRom[1586] <= 10'b0000000000;
    pxcRom[1587] <= 10'b0000000000;
    pxcRom[1588] <= 10'b0000000000;
    pxcRom[1589] <= 10'b0000000000;
    pxcRom[1590] <= 10'b0000000000;
    pxcRom[1591] <= 10'b0000000000;
    pxcRom[1592] <= 10'b0000000000;
    pxcRom[1593] <= 10'b0000000000;
    pxcRom[1594] <= 10'b0000000000;
    pxcRom[1595] <= 10'b0000000000;
    pxcRom[1596] <= 10'b0000000000;
    pxcRom[1597] <= 10'b0000000000;
    pxcRom[1598] <= 10'b0000000000;
    pxcRom[1599] <= 10'b0000000000;
    pxcRom[1600] <= 10'b0000000000;
    pxcRom[1601] <= 10'b0000000000;
    pxcRom[1602] <= 10'b0000000000;
    pxcRom[1603] <= 10'b0000000000;
    pxcRom[1604] <= 10'b0000000000;
    pxcRom[1605] <= 10'b0000000000;
    pxcRom[1606] <= 10'b0000000000;
    pxcRom[1607] <= 10'b0000000000;
    pxcRom[1608] <= 10'b0000000000;
    pxcRom[1609] <= 10'b0000000000;
    pxcRom[1610] <= 10'b0000000000;
    pxcRom[1611] <= 10'b0000000000;
    pxcRom[1612] <= 10'b0000000000;
    pxcRom[1613] <= 10'b0000000000;
    pxcRom[1614] <= 10'b0000000000;
    pxcRom[1615] <= 10'b0000000000;
    pxcRom[1616] <= 10'b0000000000;
    pxcRom[1617] <= 10'b0000000000;
    pxcRom[1618] <= 10'b0000000000;
    pxcRom[1619] <= 10'b0000000000;
    pxcRom[1620] <= 10'b0000000000;
    pxcRom[1621] <= 10'b0000000000;
    pxcRom[1622] <= 10'b0000000000;
    pxcRom[1623] <= 10'b0000000000;
    pxcRom[1624] <= 10'b0000000000;
    pxcRom[1625] <= 10'b0000000000;
    pxcRom[1626] <= 10'b0000000000;
    pxcRom[1627] <= 10'b0000000000;
    pxcRom[1628] <= 10'b0000000000;
    pxcRom[1629] <= 10'b0000000000;
    pxcRom[1630] <= 10'b0000000000;
    pxcRom[1631] <= 10'b0000000000;
    pxcRom[1632] <= 10'b0000000000;
    pxcRom[1633] <= 10'b0000000000;
    pxcRom[1634] <= 10'b0000000000;
    pxcRom[1635] <= 10'b0000000001;
    pxcRom[1636] <= 10'b0000000001;
    pxcRom[1637] <= 10'b0000000001;
    pxcRom[1638] <= 10'b0000000001;
    pxcRom[1639] <= 10'b0000000001;
    pxcRom[1640] <= 10'b0000000001;
    pxcRom[1641] <= 10'b0000000000;
    pxcRom[1642] <= 10'b0000000000;
    pxcRom[1643] <= 10'b0000000000;
    pxcRom[1644] <= 10'b0000000000;
    pxcRom[1645] <= 10'b0000000000;
    pxcRom[1646] <= 10'b0000000000;
    pxcRom[1647] <= 10'b0000000000;
    pxcRom[1648] <= 10'b0000000000;
    pxcRom[1649] <= 10'b0000000000;
    pxcRom[1650] <= 10'b0000000000;
    pxcRom[1651] <= 10'b0000000000;
    pxcRom[1652] <= 10'b0000000000;
    pxcRom[1653] <= 10'b0000000000;
    pxcRom[1654] <= 10'b0000000000;
    pxcRom[1655] <= 10'b0000000000;
    pxcRom[1656] <= 10'b0000000000;
    pxcRom[1657] <= 10'b0000000000;
    pxcRom[1658] <= 10'b0000000000;
    pxcRom[1659] <= 10'b0000000001;
    pxcRom[1660] <= 10'b0000000010;
    pxcRom[1661] <= 10'b0000000100;
    pxcRom[1662] <= 10'b0000000111;
    pxcRom[1663] <= 10'b0000001010;
    pxcRom[1664] <= 10'b0000001101;
    pxcRom[1665] <= 10'b0000001111;
    pxcRom[1666] <= 10'b0000010001;
    pxcRom[1667] <= 10'b0000010000;
    pxcRom[1668] <= 10'b0000001110;
    pxcRom[1669] <= 10'b0000001011;
    pxcRom[1670] <= 10'b0000000111;
    pxcRom[1671] <= 10'b0000000100;
    pxcRom[1672] <= 10'b0000000010;
    pxcRom[1673] <= 10'b0000000001;
    pxcRom[1674] <= 10'b0000000000;
    pxcRom[1675] <= 10'b0000000000;
    pxcRom[1676] <= 10'b0000000000;
    pxcRom[1677] <= 10'b0000000000;
    pxcRom[1678] <= 10'b0000000000;
    pxcRom[1679] <= 10'b0000000000;
    pxcRom[1680] <= 10'b0000000000;
    pxcRom[1681] <= 10'b0000000000;
    pxcRom[1682] <= 10'b0000000000;
    pxcRom[1683] <= 10'b0000000000;
    pxcRom[1684] <= 10'b0000000000;
    pxcRom[1685] <= 10'b0000000000;
    pxcRom[1686] <= 10'b0000000010;
    pxcRom[1687] <= 10'b0000000100;
    pxcRom[1688] <= 10'b0000001000;
    pxcRom[1689] <= 10'b0000001111;
    pxcRom[1690] <= 10'b0000010110;
    pxcRom[1691] <= 10'b0000100000;
    pxcRom[1692] <= 10'b0000101011;
    pxcRom[1693] <= 10'b0000110101;
    pxcRom[1694] <= 10'b0000111001;
    pxcRom[1695] <= 10'b0000111000;
    pxcRom[1696] <= 10'b0000110001;
    pxcRom[1697] <= 10'b0000100110;
    pxcRom[1698] <= 10'b0000011010;
    pxcRom[1699] <= 10'b0000010000;
    pxcRom[1700] <= 10'b0000001001;
    pxcRom[1701] <= 10'b0000000100;
    pxcRom[1702] <= 10'b0000000001;
    pxcRom[1703] <= 10'b0000000000;
    pxcRom[1704] <= 10'b0000000000;
    pxcRom[1705] <= 10'b0000000000;
    pxcRom[1706] <= 10'b0000000000;
    pxcRom[1707] <= 10'b0000000000;
    pxcRom[1708] <= 10'b0000000000;
    pxcRom[1709] <= 10'b0000000000;
    pxcRom[1710] <= 10'b0000000000;
    pxcRom[1711] <= 10'b0000000000;
    pxcRom[1712] <= 10'b0000000000;
    pxcRom[1713] <= 10'b0000000001;
    pxcRom[1714] <= 10'b0000000100;
    pxcRom[1715] <= 10'b0000001001;
    pxcRom[1716] <= 10'b0000010001;
    pxcRom[1717] <= 10'b0000011011;
    pxcRom[1718] <= 10'b0000101000;
    pxcRom[1719] <= 10'b0000111000;
    pxcRom[1720] <= 10'b0001000110;
    pxcRom[1721] <= 10'b0001010100;
    pxcRom[1722] <= 10'b0001011100;
    pxcRom[1723] <= 10'b0001011110;
    pxcRom[1724] <= 10'b0001010100;
    pxcRom[1725] <= 10'b0001000010;
    pxcRom[1726] <= 10'b0000101110;
    pxcRom[1727] <= 10'b0000011101;
    pxcRom[1728] <= 10'b0000010001;
    pxcRom[1729] <= 10'b0000001001;
    pxcRom[1730] <= 10'b0000000011;
    pxcRom[1731] <= 10'b0000000000;
    pxcRom[1732] <= 10'b0000000000;
    pxcRom[1733] <= 10'b0000000000;
    pxcRom[1734] <= 10'b0000000000;
    pxcRom[1735] <= 10'b0000000000;
    pxcRom[1736] <= 10'b0000000000;
    pxcRom[1737] <= 10'b0000000000;
    pxcRom[1738] <= 10'b0000000000;
    pxcRom[1739] <= 10'b0000000000;
    pxcRom[1740] <= 10'b0000000000;
    pxcRom[1741] <= 10'b0000000010;
    pxcRom[1742] <= 10'b0000001000;
    pxcRom[1743] <= 10'b0000001111;
    pxcRom[1744] <= 10'b0000011001;
    pxcRom[1745] <= 10'b0000100101;
    pxcRom[1746] <= 10'b0000110011;
    pxcRom[1747] <= 10'b0001000001;
    pxcRom[1748] <= 10'b0001001101;
    pxcRom[1749] <= 10'b0001010101;
    pxcRom[1750] <= 10'b0001011011;
    pxcRom[1751] <= 10'b0001011101;
    pxcRom[1752] <= 10'b0001011100;
    pxcRom[1753] <= 10'b0001010000;
    pxcRom[1754] <= 10'b0000111101;
    pxcRom[1755] <= 10'b0000101001;
    pxcRom[1756] <= 10'b0000011000;
    pxcRom[1757] <= 10'b0000001101;
    pxcRom[1758] <= 10'b0000000101;
    pxcRom[1759] <= 10'b0000000001;
    pxcRom[1760] <= 10'b0000000000;
    pxcRom[1761] <= 10'b0000000000;
    pxcRom[1762] <= 10'b0000000000;
    pxcRom[1763] <= 10'b0000000000;
    pxcRom[1764] <= 10'b0000000000;
    pxcRom[1765] <= 10'b0000000000;
    pxcRom[1766] <= 10'b0000000000;
    pxcRom[1767] <= 10'b0000000000;
    pxcRom[1768] <= 10'b0000000001;
    pxcRom[1769] <= 10'b0000000100;
    pxcRom[1770] <= 10'b0000001010;
    pxcRom[1771] <= 10'b0000010001;
    pxcRom[1772] <= 10'b0000011011;
    pxcRom[1773] <= 10'b0000100101;
    pxcRom[1774] <= 10'b0000101111;
    pxcRom[1775] <= 10'b0000110111;
    pxcRom[1776] <= 10'b0000111010;
    pxcRom[1777] <= 10'b0000111010;
    pxcRom[1778] <= 10'b0000111100;
    pxcRom[1779] <= 10'b0001000000;
    pxcRom[1780] <= 10'b0001000110;
    pxcRom[1781] <= 10'b0001001010;
    pxcRom[1782] <= 10'b0001000001;
    pxcRom[1783] <= 10'b0000110001;
    pxcRom[1784] <= 10'b0000011110;
    pxcRom[1785] <= 10'b0000010001;
    pxcRom[1786] <= 10'b0000000111;
    pxcRom[1787] <= 10'b0000000010;
    pxcRom[1788] <= 10'b0000000000;
    pxcRom[1789] <= 10'b0000000000;
    pxcRom[1790] <= 10'b0000000000;
    pxcRom[1791] <= 10'b0000000000;
    pxcRom[1792] <= 10'b0000000000;
    pxcRom[1793] <= 10'b0000000000;
    pxcRom[1794] <= 10'b0000000000;
    pxcRom[1795] <= 10'b0000000000;
    pxcRom[1796] <= 10'b0000000001;
    pxcRom[1797] <= 10'b0000000100;
    pxcRom[1798] <= 10'b0000001001;
    pxcRom[1799] <= 10'b0000010000;
    pxcRom[1800] <= 10'b0000010111;
    pxcRom[1801] <= 10'b0000011101;
    pxcRom[1802] <= 10'b0000100011;
    pxcRom[1803] <= 10'b0000100100;
    pxcRom[1804] <= 10'b0000100100;
    pxcRom[1805] <= 10'b0000100011;
    pxcRom[1806] <= 10'b0000100100;
    pxcRom[1807] <= 10'b0000101001;
    pxcRom[1808] <= 10'b0000110011;
    pxcRom[1809] <= 10'b0000111111;
    pxcRom[1810] <= 10'b0001000001;
    pxcRom[1811] <= 10'b0000110101;
    pxcRom[1812] <= 10'b0000100010;
    pxcRom[1813] <= 10'b0000010011;
    pxcRom[1814] <= 10'b0000001000;
    pxcRom[1815] <= 10'b0000000010;
    pxcRom[1816] <= 10'b0000000000;
    pxcRom[1817] <= 10'b0000000000;
    pxcRom[1818] <= 10'b0000000000;
    pxcRom[1819] <= 10'b0000000000;
    pxcRom[1820] <= 10'b0000000000;
    pxcRom[1821] <= 10'b0000000000;
    pxcRom[1822] <= 10'b0000000000;
    pxcRom[1823] <= 10'b0000000000;
    pxcRom[1824] <= 10'b0000000001;
    pxcRom[1825] <= 10'b0000000011;
    pxcRom[1826] <= 10'b0000001000;
    pxcRom[1827] <= 10'b0000001100;
    pxcRom[1828] <= 10'b0000010000;
    pxcRom[1829] <= 10'b0000010011;
    pxcRom[1830] <= 10'b0000010110;
    pxcRom[1831] <= 10'b0000010101;
    pxcRom[1832] <= 10'b0000010100;
    pxcRom[1833] <= 10'b0000010011;
    pxcRom[1834] <= 10'b0000010101;
    pxcRom[1835] <= 10'b0000011101;
    pxcRom[1836] <= 10'b0000101010;
    pxcRom[1837] <= 10'b0000111011;
    pxcRom[1838] <= 10'b0001000010;
    pxcRom[1839] <= 10'b0000110111;
    pxcRom[1840] <= 10'b0000100011;
    pxcRom[1841] <= 10'b0000010010;
    pxcRom[1842] <= 10'b0000001000;
    pxcRom[1843] <= 10'b0000000010;
    pxcRom[1844] <= 10'b0000000000;
    pxcRom[1845] <= 10'b0000000000;
    pxcRom[1846] <= 10'b0000000000;
    pxcRom[1847] <= 10'b0000000000;
    pxcRom[1848] <= 10'b0000000000;
    pxcRom[1849] <= 10'b0000000000;
    pxcRom[1850] <= 10'b0000000000;
    pxcRom[1851] <= 10'b0000000000;
    pxcRom[1852] <= 10'b0000000000;
    pxcRom[1853] <= 10'b0000000011;
    pxcRom[1854] <= 10'b0000000101;
    pxcRom[1855] <= 10'b0000001000;
    pxcRom[1856] <= 10'b0000001010;
    pxcRom[1857] <= 10'b0000001011;
    pxcRom[1858] <= 10'b0000001100;
    pxcRom[1859] <= 10'b0000001011;
    pxcRom[1860] <= 10'b0000001010;
    pxcRom[1861] <= 10'b0000001010;
    pxcRom[1862] <= 10'b0000001111;
    pxcRom[1863] <= 10'b0000011000;
    pxcRom[1864] <= 10'b0000101001;
    pxcRom[1865] <= 10'b0000111100;
    pxcRom[1866] <= 10'b0001000010;
    pxcRom[1867] <= 10'b0000110110;
    pxcRom[1868] <= 10'b0000100010;
    pxcRom[1869] <= 10'b0000010001;
    pxcRom[1870] <= 10'b0000000111;
    pxcRom[1871] <= 10'b0000000010;
    pxcRom[1872] <= 10'b0000000000;
    pxcRom[1873] <= 10'b0000000000;
    pxcRom[1874] <= 10'b0000000000;
    pxcRom[1875] <= 10'b0000000000;
    pxcRom[1876] <= 10'b0000000000;
    pxcRom[1877] <= 10'b0000000000;
    pxcRom[1878] <= 10'b0000000000;
    pxcRom[1879] <= 10'b0000000000;
    pxcRom[1880] <= 10'b0000000000;
    pxcRom[1881] <= 10'b0000000001;
    pxcRom[1882] <= 10'b0000000011;
    pxcRom[1883] <= 10'b0000000100;
    pxcRom[1884] <= 10'b0000000101;
    pxcRom[1885] <= 10'b0000000110;
    pxcRom[1886] <= 10'b0000000110;
    pxcRom[1887] <= 10'b0000000110;
    pxcRom[1888] <= 10'b0000000110;
    pxcRom[1889] <= 10'b0000001000;
    pxcRom[1890] <= 10'b0000001111;
    pxcRom[1891] <= 10'b0000011011;
    pxcRom[1892] <= 10'b0000101101;
    pxcRom[1893] <= 10'b0000111111;
    pxcRom[1894] <= 10'b0001000011;
    pxcRom[1895] <= 10'b0000110011;
    pxcRom[1896] <= 10'b0000011110;
    pxcRom[1897] <= 10'b0000001111;
    pxcRom[1898] <= 10'b0000000110;
    pxcRom[1899] <= 10'b0000000001;
    pxcRom[1900] <= 10'b0000000000;
    pxcRom[1901] <= 10'b0000000000;
    pxcRom[1902] <= 10'b0000000000;
    pxcRom[1903] <= 10'b0000000000;
    pxcRom[1904] <= 10'b0000000000;
    pxcRom[1905] <= 10'b0000000000;
    pxcRom[1906] <= 10'b0000000000;
    pxcRom[1907] <= 10'b0000000000;
    pxcRom[1908] <= 10'b0000000000;
    pxcRom[1909] <= 10'b0000000001;
    pxcRom[1910] <= 10'b0000000001;
    pxcRom[1911] <= 10'b0000000010;
    pxcRom[1912] <= 10'b0000000011;
    pxcRom[1913] <= 10'b0000000100;
    pxcRom[1914] <= 10'b0000000101;
    pxcRom[1915] <= 10'b0000000110;
    pxcRom[1916] <= 10'b0000000111;
    pxcRom[1917] <= 10'b0000001100;
    pxcRom[1918] <= 10'b0000010101;
    pxcRom[1919] <= 10'b0000100011;
    pxcRom[1920] <= 10'b0000110101;
    pxcRom[1921] <= 10'b0001000100;
    pxcRom[1922] <= 10'b0001000001;
    pxcRom[1923] <= 10'b0000101110;
    pxcRom[1924] <= 10'b0000011010;
    pxcRom[1925] <= 10'b0000001100;
    pxcRom[1926] <= 10'b0000000100;
    pxcRom[1927] <= 10'b0000000001;
    pxcRom[1928] <= 10'b0000000000;
    pxcRom[1929] <= 10'b0000000000;
    pxcRom[1930] <= 10'b0000000000;
    pxcRom[1931] <= 10'b0000000000;
    pxcRom[1932] <= 10'b0000000000;
    pxcRom[1933] <= 10'b0000000000;
    pxcRom[1934] <= 10'b0000000000;
    pxcRom[1935] <= 10'b0000000000;
    pxcRom[1936] <= 10'b0000000000;
    pxcRom[1937] <= 10'b0000000000;
    pxcRom[1938] <= 10'b0000000001;
    pxcRom[1939] <= 10'b0000000011;
    pxcRom[1940] <= 10'b0000000100;
    pxcRom[1941] <= 10'b0000000110;
    pxcRom[1942] <= 10'b0000001001;
    pxcRom[1943] <= 10'b0000001100;
    pxcRom[1944] <= 10'b0000010001;
    pxcRom[1945] <= 10'b0000011000;
    pxcRom[1946] <= 10'b0000100010;
    pxcRom[1947] <= 10'b0000110000;
    pxcRom[1948] <= 10'b0001000000;
    pxcRom[1949] <= 10'b0001000111;
    pxcRom[1950] <= 10'b0000111001;
    pxcRom[1951] <= 10'b0000100110;
    pxcRom[1952] <= 10'b0000010101;
    pxcRom[1953] <= 10'b0000001001;
    pxcRom[1954] <= 10'b0000000011;
    pxcRom[1955] <= 10'b0000000001;
    pxcRom[1956] <= 10'b0000000001;
    pxcRom[1957] <= 10'b0000000000;
    pxcRom[1958] <= 10'b0000000000;
    pxcRom[1959] <= 10'b0000000000;
    pxcRom[1960] <= 10'b0000000000;
    pxcRom[1961] <= 10'b0000000000;
    pxcRom[1962] <= 10'b0000000000;
    pxcRom[1963] <= 10'b0000000000;
    pxcRom[1964] <= 10'b0000000000;
    pxcRom[1965] <= 10'b0000000001;
    pxcRom[1966] <= 10'b0000000011;
    pxcRom[1967] <= 10'b0000000111;
    pxcRom[1968] <= 10'b0000001011;
    pxcRom[1969] <= 10'b0000010000;
    pxcRom[1970] <= 10'b0000010101;
    pxcRom[1971] <= 10'b0000011101;
    pxcRom[1972] <= 10'b0000100101;
    pxcRom[1973] <= 10'b0000101111;
    pxcRom[1974] <= 10'b0000111010;
    pxcRom[1975] <= 10'b0001000110;
    pxcRom[1976] <= 10'b0001001100;
    pxcRom[1977] <= 10'b0001000101;
    pxcRom[1978] <= 10'b0000110011;
    pxcRom[1979] <= 10'b0000100000;
    pxcRom[1980] <= 10'b0000010001;
    pxcRom[1981] <= 10'b0000001000;
    pxcRom[1982] <= 10'b0000000100;
    pxcRom[1983] <= 10'b0000000010;
    pxcRom[1984] <= 10'b0000000001;
    pxcRom[1985] <= 10'b0000000001;
    pxcRom[1986] <= 10'b0000000000;
    pxcRom[1987] <= 10'b0000000000;
    pxcRom[1988] <= 10'b0000000000;
    pxcRom[1989] <= 10'b0000000000;
    pxcRom[1990] <= 10'b0000000000;
    pxcRom[1991] <= 10'b0000000000;
    pxcRom[1992] <= 10'b0000000001;
    pxcRom[1993] <= 10'b0000000100;
    pxcRom[1994] <= 10'b0000001001;
    pxcRom[1995] <= 10'b0000010000;
    pxcRom[1996] <= 10'b0000010111;
    pxcRom[1997] <= 10'b0000100000;
    pxcRom[1998] <= 10'b0000101010;
    pxcRom[1999] <= 10'b0000110101;
    pxcRom[2000] <= 10'b0001000011;
    pxcRom[2001] <= 10'b0001010001;
    pxcRom[2002] <= 10'b0001011011;
    pxcRom[2003] <= 10'b0001011101;
    pxcRom[2004] <= 10'b0001010010;
    pxcRom[2005] <= 10'b0001000001;
    pxcRom[2006] <= 10'b0000101101;
    pxcRom[2007] <= 10'b0000011100;
    pxcRom[2008] <= 10'b0000010000;
    pxcRom[2009] <= 10'b0000001001;
    pxcRom[2010] <= 10'b0000000110;
    pxcRom[2011] <= 10'b0000000100;
    pxcRom[2012] <= 10'b0000000011;
    pxcRom[2013] <= 10'b0000000001;
    pxcRom[2014] <= 10'b0000000000;
    pxcRom[2015] <= 10'b0000000000;
    pxcRom[2016] <= 10'b0000000000;
    pxcRom[2017] <= 10'b0000000000;
    pxcRom[2018] <= 10'b0000000000;
    pxcRom[2019] <= 10'b0000000000;
    pxcRom[2020] <= 10'b0000000011;
    pxcRom[2021] <= 10'b0000001001;
    pxcRom[2022] <= 10'b0000010001;
    pxcRom[2023] <= 10'b0000011100;
    pxcRom[2024] <= 10'b0000101000;
    pxcRom[2025] <= 10'b0000110100;
    pxcRom[2026] <= 10'b0001000000;
    pxcRom[2027] <= 10'b0001001110;
    pxcRom[2028] <= 10'b0001011110;
    pxcRom[2029] <= 10'b0001101001;
    pxcRom[2030] <= 10'b0001101100;
    pxcRom[2031] <= 10'b0001100001;
    pxcRom[2032] <= 10'b0001001111;
    pxcRom[2033] <= 10'b0000111100;
    pxcRom[2034] <= 10'b0000101011;
    pxcRom[2035] <= 10'b0000011101;
    pxcRom[2036] <= 10'b0000010100;
    pxcRom[2037] <= 10'b0000001110;
    pxcRom[2038] <= 10'b0000001010;
    pxcRom[2039] <= 10'b0000001000;
    pxcRom[2040] <= 10'b0000000101;
    pxcRom[2041] <= 10'b0000000010;
    pxcRom[2042] <= 10'b0000000000;
    pxcRom[2043] <= 10'b0000000000;
    pxcRom[2044] <= 10'b0000000000;
    pxcRom[2045] <= 10'b0000000000;
    pxcRom[2046] <= 10'b0000000000;
    pxcRom[2047] <= 10'b0000000001;
    pxcRom[2048] <= 10'b0000000110;
    pxcRom[2049] <= 10'b0000001111;
    pxcRom[2050] <= 10'b0000011011;
    pxcRom[2051] <= 10'b0000101010;
    pxcRom[2052] <= 10'b0000110101;
    pxcRom[2053] <= 10'b0001000000;
    pxcRom[2054] <= 10'b0001001011;
    pxcRom[2055] <= 10'b0001011000;
    pxcRom[2056] <= 10'b0001100001;
    pxcRom[2057] <= 10'b0001101001;
    pxcRom[2058] <= 10'b0001100110;
    pxcRom[2059] <= 10'b0001011010;
    pxcRom[2060] <= 10'b0001001100;
    pxcRom[2061] <= 10'b0000111101;
    pxcRom[2062] <= 10'b0000110000;
    pxcRom[2063] <= 10'b0000100100;
    pxcRom[2064] <= 10'b0000011100;
    pxcRom[2065] <= 10'b0000010110;
    pxcRom[2066] <= 10'b0000010001;
    pxcRom[2067] <= 10'b0000001100;
    pxcRom[2068] <= 10'b0000001000;
    pxcRom[2069] <= 10'b0000000100;
    pxcRom[2070] <= 10'b0000000000;
    pxcRom[2071] <= 10'b0000000000;
    pxcRom[2072] <= 10'b0000000000;
    pxcRom[2073] <= 10'b0000000000;
    pxcRom[2074] <= 10'b0000000000;
    pxcRom[2075] <= 10'b0000000010;
    pxcRom[2076] <= 10'b0000001001;
    pxcRom[2077] <= 10'b0000010100;
    pxcRom[2078] <= 10'b0000100100;
    pxcRom[2079] <= 10'b0000110011;
    pxcRom[2080] <= 10'b0001000000;
    pxcRom[2081] <= 10'b0001001010;
    pxcRom[2082] <= 10'b0001010001;
    pxcRom[2083] <= 10'b0001011001;
    pxcRom[2084] <= 10'b0001100001;
    pxcRom[2085] <= 10'b0001100011;
    pxcRom[2086] <= 10'b0001011101;
    pxcRom[2087] <= 10'b0001010100;
    pxcRom[2088] <= 10'b0001001011;
    pxcRom[2089] <= 10'b0001000010;
    pxcRom[2090] <= 10'b0000111000;
    pxcRom[2091] <= 10'b0000101111;
    pxcRom[2092] <= 10'b0000100111;
    pxcRom[2093] <= 10'b0000100000;
    pxcRom[2094] <= 10'b0000011001;
    pxcRom[2095] <= 10'b0000010010;
    pxcRom[2096] <= 10'b0000001011;
    pxcRom[2097] <= 10'b0000000100;
    pxcRom[2098] <= 10'b0000000000;
    pxcRom[2099] <= 10'b0000000000;
    pxcRom[2100] <= 10'b0000000000;
    pxcRom[2101] <= 10'b0000000000;
    pxcRom[2102] <= 10'b0000000000;
    pxcRom[2103] <= 10'b0000000011;
    pxcRom[2104] <= 10'b0000001011;
    pxcRom[2105] <= 10'b0000010111;
    pxcRom[2106] <= 10'b0000101001;
    pxcRom[2107] <= 10'b0000111100;
    pxcRom[2108] <= 10'b0001001101;
    pxcRom[2109] <= 10'b0001011001;
    pxcRom[2110] <= 10'b0001100001;
    pxcRom[2111] <= 10'b0001100101;
    pxcRom[2112] <= 10'b0001100100;
    pxcRom[2113] <= 10'b0001100000;
    pxcRom[2114] <= 10'b0001010111;
    pxcRom[2115] <= 10'b0001001101;
    pxcRom[2116] <= 10'b0001000111;
    pxcRom[2117] <= 10'b0001000010;
    pxcRom[2118] <= 10'b0000111101;
    pxcRom[2119] <= 10'b0000111000;
    pxcRom[2120] <= 10'b0000101111;
    pxcRom[2121] <= 10'b0000100111;
    pxcRom[2122] <= 10'b0000011101;
    pxcRom[2123] <= 10'b0000010100;
    pxcRom[2124] <= 10'b0000001011;
    pxcRom[2125] <= 10'b0000000100;
    pxcRom[2126] <= 10'b0000000000;
    pxcRom[2127] <= 10'b0000000000;
    pxcRom[2128] <= 10'b0000000000;
    pxcRom[2129] <= 10'b0000000000;
    pxcRom[2130] <= 10'b0000000000;
    pxcRom[2131] <= 10'b0000000011;
    pxcRom[2132] <= 10'b0000001011;
    pxcRom[2133] <= 10'b0000010111;
    pxcRom[2134] <= 10'b0000101001;
    pxcRom[2135] <= 10'b0000111110;
    pxcRom[2136] <= 10'b0001010101;
    pxcRom[2137] <= 10'b0001100101;
    pxcRom[2138] <= 10'b0001101010;
    pxcRom[2139] <= 10'b0001101001;
    pxcRom[2140] <= 10'b0001011111;
    pxcRom[2141] <= 10'b0001010000;
    pxcRom[2142] <= 10'b0001000100;
    pxcRom[2143] <= 10'b0000111100;
    pxcRom[2144] <= 10'b0000111001;
    pxcRom[2145] <= 10'b0000110111;
    pxcRom[2146] <= 10'b0000110111;
    pxcRom[2147] <= 10'b0000110011;
    pxcRom[2148] <= 10'b0000101110;
    pxcRom[2149] <= 10'b0000100100;
    pxcRom[2150] <= 10'b0000011011;
    pxcRom[2151] <= 10'b0000010001;
    pxcRom[2152] <= 10'b0000001001;
    pxcRom[2153] <= 10'b0000000011;
    pxcRom[2154] <= 10'b0000000000;
    pxcRom[2155] <= 10'b0000000000;
    pxcRom[2156] <= 10'b0000000000;
    pxcRom[2157] <= 10'b0000000000;
    pxcRom[2158] <= 10'b0000000000;
    pxcRom[2159] <= 10'b0000000010;
    pxcRom[2160] <= 10'b0000001001;
    pxcRom[2161] <= 10'b0000010010;
    pxcRom[2162] <= 10'b0000100001;
    pxcRom[2163] <= 10'b0000110011;
    pxcRom[2164] <= 10'b0001000111;
    pxcRom[2165] <= 10'b0001010101;
    pxcRom[2166] <= 10'b0001010111;
    pxcRom[2167] <= 10'b0001010000;
    pxcRom[2168] <= 10'b0001000100;
    pxcRom[2169] <= 10'b0000110111;
    pxcRom[2170] <= 10'b0000101101;
    pxcRom[2171] <= 10'b0000100111;
    pxcRom[2172] <= 10'b0000100101;
    pxcRom[2173] <= 10'b0000100110;
    pxcRom[2174] <= 10'b0000100111;
    pxcRom[2175] <= 10'b0000100110;
    pxcRom[2176] <= 10'b0000100010;
    pxcRom[2177] <= 10'b0000011010;
    pxcRom[2178] <= 10'b0000010010;
    pxcRom[2179] <= 10'b0000001100;
    pxcRom[2180] <= 10'b0000000110;
    pxcRom[2181] <= 10'b0000000001;
    pxcRom[2182] <= 10'b0000000000;
    pxcRom[2183] <= 10'b0000000000;
    pxcRom[2184] <= 10'b0000000000;
    pxcRom[2185] <= 10'b0000000000;
    pxcRom[2186] <= 10'b0000000000;
    pxcRom[2187] <= 10'b0000000001;
    pxcRom[2188] <= 10'b0000000101;
    pxcRom[2189] <= 10'b0000001011;
    pxcRom[2190] <= 10'b0000010100;
    pxcRom[2191] <= 10'b0000100000;
    pxcRom[2192] <= 10'b0000101011;
    pxcRom[2193] <= 10'b0000110001;
    pxcRom[2194] <= 10'b0000110010;
    pxcRom[2195] <= 10'b0000101101;
    pxcRom[2196] <= 10'b0000100101;
    pxcRom[2197] <= 10'b0000011110;
    pxcRom[2198] <= 10'b0000011000;
    pxcRom[2199] <= 10'b0000010101;
    pxcRom[2200] <= 10'b0000010100;
    pxcRom[2201] <= 10'b0000010101;
    pxcRom[2202] <= 10'b0000010110;
    pxcRom[2203] <= 10'b0000010101;
    pxcRom[2204] <= 10'b0000010011;
    pxcRom[2205] <= 10'b0000001110;
    pxcRom[2206] <= 10'b0000001010;
    pxcRom[2207] <= 10'b0000000110;
    pxcRom[2208] <= 10'b0000000011;
    pxcRom[2209] <= 10'b0000000000;
    pxcRom[2210] <= 10'b0000000000;
    pxcRom[2211] <= 10'b0000000000;
    pxcRom[2212] <= 10'b0000000000;
    pxcRom[2213] <= 10'b0000000000;
    pxcRom[2214] <= 10'b0000000000;
    pxcRom[2215] <= 10'b0000000000;
    pxcRom[2216] <= 10'b0000000001;
    pxcRom[2217] <= 10'b0000000011;
    pxcRom[2218] <= 10'b0000000110;
    pxcRom[2219] <= 10'b0000001010;
    pxcRom[2220] <= 10'b0000001110;
    pxcRom[2221] <= 10'b0000010000;
    pxcRom[2222] <= 10'b0000010000;
    pxcRom[2223] <= 10'b0000001111;
    pxcRom[2224] <= 10'b0000001101;
    pxcRom[2225] <= 10'b0000001011;
    pxcRom[2226] <= 10'b0000001001;
    pxcRom[2227] <= 10'b0000001000;
    pxcRom[2228] <= 10'b0000001000;
    pxcRom[2229] <= 10'b0000001000;
    pxcRom[2230] <= 10'b0000001000;
    pxcRom[2231] <= 10'b0000000111;
    pxcRom[2232] <= 10'b0000000110;
    pxcRom[2233] <= 10'b0000000101;
    pxcRom[2234] <= 10'b0000000011;
    pxcRom[2235] <= 10'b0000000010;
    pxcRom[2236] <= 10'b0000000000;
    pxcRom[2237] <= 10'b0000000000;
    pxcRom[2238] <= 10'b0000000000;
    pxcRom[2239] <= 10'b0000000000;
    pxcRom[2240] <= 10'b0000000000;
    pxcRom[2241] <= 10'b0000000000;
    pxcRom[2242] <= 10'b0000000000;
    pxcRom[2243] <= 10'b0000000000;
    pxcRom[2244] <= 10'b0000000000;
    pxcRom[2245] <= 10'b0000000000;
    pxcRom[2246] <= 10'b0000000000;
    pxcRom[2247] <= 10'b0000000000;
    pxcRom[2248] <= 10'b0000000001;
    pxcRom[2249] <= 10'b0000000001;
    pxcRom[2250] <= 10'b0000000001;
    pxcRom[2251] <= 10'b0000000001;
    pxcRom[2252] <= 10'b0000000001;
    pxcRom[2253] <= 10'b0000000001;
    pxcRom[2254] <= 10'b0000000001;
    pxcRom[2255] <= 10'b0000000001;
    pxcRom[2256] <= 10'b0000000001;
    pxcRom[2257] <= 10'b0000000001;
    pxcRom[2258] <= 10'b0000000001;
    pxcRom[2259] <= 10'b0000000001;
    pxcRom[2260] <= 10'b0000000000;
    pxcRom[2261] <= 10'b0000000000;
    pxcRom[2262] <= 10'b0000000000;
    pxcRom[2263] <= 10'b0000000000;
    pxcRom[2264] <= 10'b0000000000;
    pxcRom[2265] <= 10'b0000000000;
    pxcRom[2266] <= 10'b0000000000;
    pxcRom[2267] <= 10'b0000000000;
    pxcRom[2268] <= 10'b0000000000;
    pxcRom[2269] <= 10'b0000000000;
    pxcRom[2270] <= 10'b0000000000;
    pxcRom[2271] <= 10'b0000000000;
    pxcRom[2272] <= 10'b0000000000;
    pxcRom[2273] <= 10'b0000000000;
    pxcRom[2274] <= 10'b0000000000;
    pxcRom[2275] <= 10'b0000000000;
    pxcRom[2276] <= 10'b0000000000;
    pxcRom[2277] <= 10'b0000000000;
    pxcRom[2278] <= 10'b0000000000;
    pxcRom[2279] <= 10'b0000000000;
    pxcRom[2280] <= 10'b0000000000;
    pxcRom[2281] <= 10'b0000000000;
    pxcRom[2282] <= 10'b0000000000;
    pxcRom[2283] <= 10'b0000000000;
    pxcRom[2284] <= 10'b0000000000;
    pxcRom[2285] <= 10'b0000000000;
    pxcRom[2286] <= 10'b0000000000;
    pxcRom[2287] <= 10'b0000000000;
    pxcRom[2288] <= 10'b0000000000;
    pxcRom[2289] <= 10'b0000000000;
    pxcRom[2290] <= 10'b0000000000;
    pxcRom[2291] <= 10'b0000000000;
    pxcRom[2292] <= 10'b0000000000;
    pxcRom[2293] <= 10'b0000000000;
    pxcRom[2294] <= 10'b0000000000;
    pxcRom[2295] <= 10'b0000000000;
    pxcRom[2296] <= 10'b0000000000;
    pxcRom[2297] <= 10'b0000000000;
    pxcRom[2298] <= 10'b0000000000;
    pxcRom[2299] <= 10'b0000000000;
    pxcRom[2300] <= 10'b0000000000;
    pxcRom[2301] <= 10'b0000000000;
    pxcRom[2302] <= 10'b0000000000;
    pxcRom[2303] <= 10'b0000000000;
    pxcRom[2304] <= 10'b0000000000;
    pxcRom[2305] <= 10'b0000000000;
    pxcRom[2306] <= 10'b0000000000;
    pxcRom[2307] <= 10'b0000000000;
    pxcRom[2308] <= 10'b0000000000;
    pxcRom[2309] <= 10'b0000000000;
    pxcRom[2310] <= 10'b0000000000;
    pxcRom[2311] <= 10'b0000000000;
    pxcRom[2312] <= 10'b0000000000;
    pxcRom[2313] <= 10'b0000000000;
    pxcRom[2314] <= 10'b0000000000;
    pxcRom[2315] <= 10'b0000000000;
    pxcRom[2316] <= 10'b0000000000;
    pxcRom[2317] <= 10'b0000000000;
    pxcRom[2318] <= 10'b0000000000;
    pxcRom[2319] <= 10'b0000000000;
    pxcRom[2320] <= 10'b0000000000;
    pxcRom[2321] <= 10'b0000000000;
    pxcRom[2322] <= 10'b0000000000;
    pxcRom[2323] <= 10'b0000000000;
    pxcRom[2324] <= 10'b0000000000;
    pxcRom[2325] <= 10'b0000000000;
    pxcRom[2326] <= 10'b0000000000;
    pxcRom[2327] <= 10'b0000000000;
    pxcRom[2328] <= 10'b0000000000;
    pxcRom[2329] <= 10'b0000000000;
    pxcRom[2330] <= 10'b0000000000;
    pxcRom[2331] <= 10'b0000000000;
    pxcRom[2332] <= 10'b0000000000;
    pxcRom[2333] <= 10'b0000000000;
    pxcRom[2334] <= 10'b0000000000;
    pxcRom[2335] <= 10'b0000000000;
    pxcRom[2336] <= 10'b0000000000;
    pxcRom[2337] <= 10'b0000000000;
    pxcRom[2338] <= 10'b0000000000;
    pxcRom[2339] <= 10'b0000000000;
    pxcRom[2340] <= 10'b0000000000;
    pxcRom[2341] <= 10'b0000000000;
    pxcRom[2342] <= 10'b0000000000;
    pxcRom[2343] <= 10'b0000000000;
    pxcRom[2344] <= 10'b0000000000;
    pxcRom[2345] <= 10'b0000000000;
    pxcRom[2346] <= 10'b0000000000;
    pxcRom[2347] <= 10'b0000000000;
    pxcRom[2348] <= 10'b0000000000;
    pxcRom[2349] <= 10'b0000000000;
    pxcRom[2350] <= 10'b0000000000;
    pxcRom[2351] <= 10'b0000000000;
    pxcRom[2352] <= 10'b0000000000;
    pxcRom[2353] <= 10'b0000000000;
    pxcRom[2354] <= 10'b0000000000;
    pxcRom[2355] <= 10'b0000000000;
    pxcRom[2356] <= 10'b0000000000;
    pxcRom[2357] <= 10'b0000000000;
    pxcRom[2358] <= 10'b0000000000;
    pxcRom[2359] <= 10'b0000000000;
    pxcRom[2360] <= 10'b0000000000;
    pxcRom[2361] <= 10'b0000000000;
    pxcRom[2362] <= 10'b0000000000;
    pxcRom[2363] <= 10'b0000000000;
    pxcRom[2364] <= 10'b0000000000;
    pxcRom[2365] <= 10'b0000000000;
    pxcRom[2366] <= 10'b0000000000;
    pxcRom[2367] <= 10'b0000000000;
    pxcRom[2368] <= 10'b0000000000;
    pxcRom[2369] <= 10'b0000000000;
    pxcRom[2370] <= 10'b0000000000;
    pxcRom[2371] <= 10'b0000000000;
    pxcRom[2372] <= 10'b0000000000;
    pxcRom[2373] <= 10'b0000000000;
    pxcRom[2374] <= 10'b0000000000;
    pxcRom[2375] <= 10'b0000000000;
    pxcRom[2376] <= 10'b0000000000;
    pxcRom[2377] <= 10'b0000000000;
    pxcRom[2378] <= 10'b0000000000;
    pxcRom[2379] <= 10'b0000000000;
    pxcRom[2380] <= 10'b0000000000;
    pxcRom[2381] <= 10'b0000000000;
    pxcRom[2382] <= 10'b0000000000;
    pxcRom[2383] <= 10'b0000000000;
    pxcRom[2384] <= 10'b0000000000;
    pxcRom[2385] <= 10'b0000000000;
    pxcRom[2386] <= 10'b0000000000;
    pxcRom[2387] <= 10'b0000000000;
    pxcRom[2388] <= 10'b0000000000;
    pxcRom[2389] <= 10'b0000000000;
    pxcRom[2390] <= 10'b0000000000;
    pxcRom[2391] <= 10'b0000000000;
    pxcRom[2392] <= 10'b0000000000;
    pxcRom[2393] <= 10'b0000000000;
    pxcRom[2394] <= 10'b0000000000;
    pxcRom[2395] <= 10'b0000000000;
    pxcRom[2396] <= 10'b0000000000;
    pxcRom[2397] <= 10'b0000000000;
    pxcRom[2398] <= 10'b0000000000;
    pxcRom[2399] <= 10'b0000000000;
    pxcRom[2400] <= 10'b0000000000;
    pxcRom[2401] <= 10'b0000000000;
    pxcRom[2402] <= 10'b0000000000;
    pxcRom[2403] <= 10'b0000000000;
    pxcRom[2404] <= 10'b0000000000;
    pxcRom[2405] <= 10'b0000000000;
    pxcRom[2406] <= 10'b0000000000;
    pxcRom[2407] <= 10'b0000000000;
    pxcRom[2408] <= 10'b0000000000;
    pxcRom[2409] <= 10'b0000000000;
    pxcRom[2410] <= 10'b0000000000;
    pxcRom[2411] <= 10'b0000000000;
    pxcRom[2412] <= 10'b0000000000;
    pxcRom[2413] <= 10'b0000000000;
    pxcRom[2414] <= 10'b0000000000;
    pxcRom[2415] <= 10'b0000000000;
    pxcRom[2416] <= 10'b0000000000;
    pxcRom[2417] <= 10'b0000000000;
    pxcRom[2418] <= 10'b0000000000;
    pxcRom[2419] <= 10'b0000000000;
    pxcRom[2420] <= 10'b0000000000;
    pxcRom[2421] <= 10'b0000000000;
    pxcRom[2422] <= 10'b0000000000;
    pxcRom[2423] <= 10'b0000000000;
    pxcRom[2424] <= 10'b0000000000;
    pxcRom[2425] <= 10'b0000000000;
    pxcRom[2426] <= 10'b0000000000;
    pxcRom[2427] <= 10'b0000000000;
    pxcRom[2428] <= 10'b0000000000;
    pxcRom[2429] <= 10'b0000000000;
    pxcRom[2430] <= 10'b0000000000;
    pxcRom[2431] <= 10'b0000000000;
    pxcRom[2432] <= 10'b0000000000;
    pxcRom[2433] <= 10'b0000000000;
    pxcRom[2434] <= 10'b0000000000;
    pxcRom[2435] <= 10'b0000000000;
    pxcRom[2436] <= 10'b0000000000;
    pxcRom[2437] <= 10'b0000000000;
    pxcRom[2438] <= 10'b0000000000;
    pxcRom[2439] <= 10'b0000000000;
    pxcRom[2440] <= 10'b0000000000;
    pxcRom[2441] <= 10'b0000000000;
    pxcRom[2442] <= 10'b0000000000;
    pxcRom[2443] <= 10'b0000000000;
    pxcRom[2444] <= 10'b0000000000;
    pxcRom[2445] <= 10'b0000000000;
    pxcRom[2446] <= 10'b0000000000;
    pxcRom[2447] <= 10'b0000000001;
    pxcRom[2448] <= 10'b0000000010;
    pxcRom[2449] <= 10'b0000000010;
    pxcRom[2450] <= 10'b0000000010;
    pxcRom[2451] <= 10'b0000000010;
    pxcRom[2452] <= 10'b0000000010;
    pxcRom[2453] <= 10'b0000000001;
    pxcRom[2454] <= 10'b0000000001;
    pxcRom[2455] <= 10'b0000000000;
    pxcRom[2456] <= 10'b0000000000;
    pxcRom[2457] <= 10'b0000000000;
    pxcRom[2458] <= 10'b0000000000;
    pxcRom[2459] <= 10'b0000000000;
    pxcRom[2460] <= 10'b0000000000;
    pxcRom[2461] <= 10'b0000000000;
    pxcRom[2462] <= 10'b0000000000;
    pxcRom[2463] <= 10'b0000000000;
    pxcRom[2464] <= 10'b0000000000;
    pxcRom[2465] <= 10'b0000000000;
    pxcRom[2466] <= 10'b0000000000;
    pxcRom[2467] <= 10'b0000000000;
    pxcRom[2468] <= 10'b0000000000;
    pxcRom[2469] <= 10'b0000000000;
    pxcRom[2470] <= 10'b0000000001;
    pxcRom[2471] <= 10'b0000000011;
    pxcRom[2472] <= 10'b0000000110;
    pxcRom[2473] <= 10'b0000001001;
    pxcRom[2474] <= 10'b0000001110;
    pxcRom[2475] <= 10'b0000010011;
    pxcRom[2476] <= 10'b0000010111;
    pxcRom[2477] <= 10'b0000011010;
    pxcRom[2478] <= 10'b0000011010;
    pxcRom[2479] <= 10'b0000011001;
    pxcRom[2480] <= 10'b0000010100;
    pxcRom[2481] <= 10'b0000001111;
    pxcRom[2482] <= 10'b0000001010;
    pxcRom[2483] <= 10'b0000000110;
    pxcRom[2484] <= 10'b0000000011;
    pxcRom[2485] <= 10'b0000000001;
    pxcRom[2486] <= 10'b0000000000;
    pxcRom[2487] <= 10'b0000000000;
    pxcRom[2488] <= 10'b0000000000;
    pxcRom[2489] <= 10'b0000000000;
    pxcRom[2490] <= 10'b0000000000;
    pxcRom[2491] <= 10'b0000000000;
    pxcRom[2492] <= 10'b0000000000;
    pxcRom[2493] <= 10'b0000000000;
    pxcRom[2494] <= 10'b0000000000;
    pxcRom[2495] <= 10'b0000000000;
    pxcRom[2496] <= 10'b0000000001;
    pxcRom[2497] <= 10'b0000000011;
    pxcRom[2498] <= 10'b0000000110;
    pxcRom[2499] <= 10'b0000001100;
    pxcRom[2500] <= 10'b0000010100;
    pxcRom[2501] <= 10'b0000011111;
    pxcRom[2502] <= 10'b0000101110;
    pxcRom[2503] <= 10'b0000111110;
    pxcRom[2504] <= 10'b0001001101;
    pxcRom[2505] <= 10'b0001011010;
    pxcRom[2506] <= 10'b0001011100;
    pxcRom[2507] <= 10'b0001010100;
    pxcRom[2508] <= 10'b0001000110;
    pxcRom[2509] <= 10'b0000110011;
    pxcRom[2510] <= 10'b0000100010;
    pxcRom[2511] <= 10'b0000010101;
    pxcRom[2512] <= 10'b0000001100;
    pxcRom[2513] <= 10'b0000000101;
    pxcRom[2514] <= 10'b0000000001;
    pxcRom[2515] <= 10'b0000000000;
    pxcRom[2516] <= 10'b0000000000;
    pxcRom[2517] <= 10'b0000000000;
    pxcRom[2518] <= 10'b0000000000;
    pxcRom[2519] <= 10'b0000000000;
    pxcRom[2520] <= 10'b0000000000;
    pxcRom[2521] <= 10'b0000000000;
    pxcRom[2522] <= 10'b0000000000;
    pxcRom[2523] <= 10'b0000000000;
    pxcRom[2524] <= 10'b0000000010;
    pxcRom[2525] <= 10'b0000000110;
    pxcRom[2526] <= 10'b0000001100;
    pxcRom[2527] <= 10'b0000010101;
    pxcRom[2528] <= 10'b0000100011;
    pxcRom[2529] <= 10'b0000110100;
    pxcRom[2530] <= 10'b0001001001;
    pxcRom[2531] <= 10'b0001011100;
    pxcRom[2532] <= 10'b0001101110;
    pxcRom[2533] <= 10'b0001111100;
    pxcRom[2534] <= 10'b0010000010;
    pxcRom[2535] <= 10'b0010000100;
    pxcRom[2536] <= 10'b0001110010;
    pxcRom[2537] <= 10'b0001010110;
    pxcRom[2538] <= 10'b0000111001;
    pxcRom[2539] <= 10'b0000100100;
    pxcRom[2540] <= 10'b0000010101;
    pxcRom[2541] <= 10'b0000001011;
    pxcRom[2542] <= 10'b0000000100;
    pxcRom[2543] <= 10'b0000000000;
    pxcRom[2544] <= 10'b0000000000;
    pxcRom[2545] <= 10'b0000000000;
    pxcRom[2546] <= 10'b0000000000;
    pxcRom[2547] <= 10'b0000000000;
    pxcRom[2548] <= 10'b0000000000;
    pxcRom[2549] <= 10'b0000000000;
    pxcRom[2550] <= 10'b0000000000;
    pxcRom[2551] <= 10'b0000000001;
    pxcRom[2552] <= 10'b0000000011;
    pxcRom[2553] <= 10'b0000001000;
    pxcRom[2554] <= 10'b0000001111;
    pxcRom[2555] <= 10'b0000011001;
    pxcRom[2556] <= 10'b0000100100;
    pxcRom[2557] <= 10'b0000110011;
    pxcRom[2558] <= 10'b0000111110;
    pxcRom[2559] <= 10'b0001000111;
    pxcRom[2560] <= 10'b0001001010;
    pxcRom[2561] <= 10'b0001001101;
    pxcRom[2562] <= 10'b0001010100;
    pxcRom[2563] <= 10'b0001100001;
    pxcRom[2564] <= 10'b0001100101;
    pxcRom[2565] <= 10'b0001011011;
    pxcRom[2566] <= 10'b0001000100;
    pxcRom[2567] <= 10'b0000101101;
    pxcRom[2568] <= 10'b0000011010;
    pxcRom[2569] <= 10'b0000001110;
    pxcRom[2570] <= 10'b0000000101;
    pxcRom[2571] <= 10'b0000000001;
    pxcRom[2572] <= 10'b0000000000;
    pxcRom[2573] <= 10'b0000000000;
    pxcRom[2574] <= 10'b0000000000;
    pxcRom[2575] <= 10'b0000000000;
    pxcRom[2576] <= 10'b0000000000;
    pxcRom[2577] <= 10'b0000000000;
    pxcRom[2578] <= 10'b0000000000;
    pxcRom[2579] <= 10'b0000000001;
    pxcRom[2580] <= 10'b0000000011;
    pxcRom[2581] <= 10'b0000000111;
    pxcRom[2582] <= 10'b0000001101;
    pxcRom[2583] <= 10'b0000010100;
    pxcRom[2584] <= 10'b0000011011;
    pxcRom[2585] <= 10'b0000100001;
    pxcRom[2586] <= 10'b0000100011;
    pxcRom[2587] <= 10'b0000100100;
    pxcRom[2588] <= 10'b0000100011;
    pxcRom[2589] <= 10'b0000100101;
    pxcRom[2590] <= 10'b0000101100;
    pxcRom[2591] <= 10'b0000111011;
    pxcRom[2592] <= 10'b0001001001;
    pxcRom[2593] <= 10'b0001010000;
    pxcRom[2594] <= 10'b0001000100;
    pxcRom[2595] <= 10'b0000101111;
    pxcRom[2596] <= 10'b0000011100;
    pxcRom[2597] <= 10'b0000001110;
    pxcRom[2598] <= 10'b0000000101;
    pxcRom[2599] <= 10'b0000000001;
    pxcRom[2600] <= 10'b0000000000;
    pxcRom[2601] <= 10'b0000000000;
    pxcRom[2602] <= 10'b0000000000;
    pxcRom[2603] <= 10'b0000000000;
    pxcRom[2604] <= 10'b0000000000;
    pxcRom[2605] <= 10'b0000000000;
    pxcRom[2606] <= 10'b0000000000;
    pxcRom[2607] <= 10'b0000000001;
    pxcRom[2608] <= 10'b0000000011;
    pxcRom[2609] <= 10'b0000000101;
    pxcRom[2610] <= 10'b0000001001;
    pxcRom[2611] <= 10'b0000001100;
    pxcRom[2612] <= 10'b0000001110;
    pxcRom[2613] <= 10'b0000010000;
    pxcRom[2614] <= 10'b0000010001;
    pxcRom[2615] <= 10'b0000010001;
    pxcRom[2616] <= 10'b0000010010;
    pxcRom[2617] <= 10'b0000010111;
    pxcRom[2618] <= 10'b0000100010;
    pxcRom[2619] <= 10'b0000110100;
    pxcRom[2620] <= 10'b0001001001;
    pxcRom[2621] <= 10'b0001010000;
    pxcRom[2622] <= 10'b0001000001;
    pxcRom[2623] <= 10'b0000101010;
    pxcRom[2624] <= 10'b0000011000;
    pxcRom[2625] <= 10'b0000001011;
    pxcRom[2626] <= 10'b0000000100;
    pxcRom[2627] <= 10'b0000000000;
    pxcRom[2628] <= 10'b0000000000;
    pxcRom[2629] <= 10'b0000000000;
    pxcRom[2630] <= 10'b0000000000;
    pxcRom[2631] <= 10'b0000000000;
    pxcRom[2632] <= 10'b0000000000;
    pxcRom[2633] <= 10'b0000000000;
    pxcRom[2634] <= 10'b0000000000;
    pxcRom[2635] <= 10'b0000000000;
    pxcRom[2636] <= 10'b0000000001;
    pxcRom[2637] <= 10'b0000000010;
    pxcRom[2638] <= 10'b0000000100;
    pxcRom[2639] <= 10'b0000000101;
    pxcRom[2640] <= 10'b0000000111;
    pxcRom[2641] <= 10'b0000001000;
    pxcRom[2642] <= 10'b0000001010;
    pxcRom[2643] <= 10'b0000001110;
    pxcRom[2644] <= 10'b0000010100;
    pxcRom[2645] <= 10'b0000011111;
    pxcRom[2646] <= 10'b0000110010;
    pxcRom[2647] <= 10'b0001001001;
    pxcRom[2648] <= 10'b0001011100;
    pxcRom[2649] <= 10'b0001010011;
    pxcRom[2650] <= 10'b0000111011;
    pxcRom[2651] <= 10'b0000100010;
    pxcRom[2652] <= 10'b0000010010;
    pxcRom[2653] <= 10'b0000000111;
    pxcRom[2654] <= 10'b0000000010;
    pxcRom[2655] <= 10'b0000000000;
    pxcRom[2656] <= 10'b0000000000;
    pxcRom[2657] <= 10'b0000000000;
    pxcRom[2658] <= 10'b0000000000;
    pxcRom[2659] <= 10'b0000000000;
    pxcRom[2660] <= 10'b0000000000;
    pxcRom[2661] <= 10'b0000000000;
    pxcRom[2662] <= 10'b0000000000;
    pxcRom[2663] <= 10'b0000000000;
    pxcRom[2664] <= 10'b0000000000;
    pxcRom[2665] <= 10'b0000000001;
    pxcRom[2666] <= 10'b0000000010;
    pxcRom[2667] <= 10'b0000000011;
    pxcRom[2668] <= 10'b0000000101;
    pxcRom[2669] <= 10'b0000001000;
    pxcRom[2670] <= 10'b0000001111;
    pxcRom[2671] <= 10'b0000011011;
    pxcRom[2672] <= 10'b0000101011;
    pxcRom[2673] <= 10'b0001000001;
    pxcRom[2674] <= 10'b0001011001;
    pxcRom[2675] <= 10'b0001101101;
    pxcRom[2676] <= 10'b0001101100;
    pxcRom[2677] <= 10'b0001010000;
    pxcRom[2678] <= 10'b0000110001;
    pxcRom[2679] <= 10'b0000011001;
    pxcRom[2680] <= 10'b0000001100;
    pxcRom[2681] <= 10'b0000000100;
    pxcRom[2682] <= 10'b0000000001;
    pxcRom[2683] <= 10'b0000000000;
    pxcRom[2684] <= 10'b0000000000;
    pxcRom[2685] <= 10'b0000000000;
    pxcRom[2686] <= 10'b0000000000;
    pxcRom[2687] <= 10'b0000000000;
    pxcRom[2688] <= 10'b0000000000;
    pxcRom[2689] <= 10'b0000000000;
    pxcRom[2690] <= 10'b0000000000;
    pxcRom[2691] <= 10'b0000000000;
    pxcRom[2692] <= 10'b0000000000;
    pxcRom[2693] <= 10'b0000000000;
    pxcRom[2694] <= 10'b0000000001;
    pxcRom[2695] <= 10'b0000000011;
    pxcRom[2696] <= 10'b0000000111;
    pxcRom[2697] <= 10'b0000010000;
    pxcRom[2698] <= 10'b0000100000;
    pxcRom[2699] <= 10'b0000110110;
    pxcRom[2700] <= 10'b0001010010;
    pxcRom[2701] <= 10'b0001110001;
    pxcRom[2702] <= 10'b0010001010;
    pxcRom[2703] <= 10'b0010001101;
    pxcRom[2704] <= 10'b0001110001;
    pxcRom[2705] <= 10'b0001001111;
    pxcRom[2706] <= 10'b0000101101;
    pxcRom[2707] <= 10'b0000010111;
    pxcRom[2708] <= 10'b0000001010;
    pxcRom[2709] <= 10'b0000000011;
    pxcRom[2710] <= 10'b0000000001;
    pxcRom[2711] <= 10'b0000000000;
    pxcRom[2712] <= 10'b0000000000;
    pxcRom[2713] <= 10'b0000000000;
    pxcRom[2714] <= 10'b0000000000;
    pxcRom[2715] <= 10'b0000000000;
    pxcRom[2716] <= 10'b0000000000;
    pxcRom[2717] <= 10'b0000000000;
    pxcRom[2718] <= 10'b0000000000;
    pxcRom[2719] <= 10'b0000000000;
    pxcRom[2720] <= 10'b0000000000;
    pxcRom[2721] <= 10'b0000000000;
    pxcRom[2722] <= 10'b0000000001;
    pxcRom[2723] <= 10'b0000000100;
    pxcRom[2724] <= 10'b0000001010;
    pxcRom[2725] <= 10'b0000011000;
    pxcRom[2726] <= 10'b0000101111;
    pxcRom[2727] <= 10'b0001001101;
    pxcRom[2728] <= 10'b0001101101;
    pxcRom[2729] <= 10'b0010001000;
    pxcRom[2730] <= 10'b0010001100;
    pxcRom[2731] <= 10'b0010000010;
    pxcRom[2732] <= 10'b0001101110;
    pxcRom[2733] <= 10'b0001010010;
    pxcRom[2734] <= 10'b0000110101;
    pxcRom[2735] <= 10'b0000011110;
    pxcRom[2736] <= 10'b0000001110;
    pxcRom[2737] <= 10'b0000000101;
    pxcRom[2738] <= 10'b0000000001;
    pxcRom[2739] <= 10'b0000000000;
    pxcRom[2740] <= 10'b0000000000;
    pxcRom[2741] <= 10'b0000000000;
    pxcRom[2742] <= 10'b0000000000;
    pxcRom[2743] <= 10'b0000000000;
    pxcRom[2744] <= 10'b0000000000;
    pxcRom[2745] <= 10'b0000000000;
    pxcRom[2746] <= 10'b0000000000;
    pxcRom[2747] <= 10'b0000000000;
    pxcRom[2748] <= 10'b0000000000;
    pxcRom[2749] <= 10'b0000000000;
    pxcRom[2750] <= 10'b0000000001;
    pxcRom[2751] <= 10'b0000000101;
    pxcRom[2752] <= 10'b0000001100;
    pxcRom[2753] <= 10'b0000011010;
    pxcRom[2754] <= 10'b0000101101;
    pxcRom[2755] <= 10'b0001000100;
    pxcRom[2756] <= 10'b0001010100;
    pxcRom[2757] <= 10'b0001011100;
    pxcRom[2758] <= 10'b0001011010;
    pxcRom[2759] <= 10'b0001011001;
    pxcRom[2760] <= 10'b0001011011;
    pxcRom[2761] <= 10'b0001010101;
    pxcRom[2762] <= 10'b0001000100;
    pxcRom[2763] <= 10'b0000101011;
    pxcRom[2764] <= 10'b0000010110;
    pxcRom[2765] <= 10'b0000001001;
    pxcRom[2766] <= 10'b0000000011;
    pxcRom[2767] <= 10'b0000000000;
    pxcRom[2768] <= 10'b0000000000;
    pxcRom[2769] <= 10'b0000000000;
    pxcRom[2770] <= 10'b0000000000;
    pxcRom[2771] <= 10'b0000000000;
    pxcRom[2772] <= 10'b0000000000;
    pxcRom[2773] <= 10'b0000000000;
    pxcRom[2774] <= 10'b0000000000;
    pxcRom[2775] <= 10'b0000000000;
    pxcRom[2776] <= 10'b0000000000;
    pxcRom[2777] <= 10'b0000000001;
    pxcRom[2778] <= 10'b0000000010;
    pxcRom[2779] <= 10'b0000000100;
    pxcRom[2780] <= 10'b0000001001;
    pxcRom[2781] <= 10'b0000010011;
    pxcRom[2782] <= 10'b0000011110;
    pxcRom[2783] <= 10'b0000100111;
    pxcRom[2784] <= 10'b0000101100;
    pxcRom[2785] <= 10'b0000101101;
    pxcRom[2786] <= 10'b0000101101;
    pxcRom[2787] <= 10'b0000110010;
    pxcRom[2788] <= 10'b0000111100;
    pxcRom[2789] <= 10'b0001001011;
    pxcRom[2790] <= 10'b0001001100;
    pxcRom[2791] <= 10'b0000111001;
    pxcRom[2792] <= 10'b0000100001;
    pxcRom[2793] <= 10'b0000001111;
    pxcRom[2794] <= 10'b0000000110;
    pxcRom[2795] <= 10'b0000000001;
    pxcRom[2796] <= 10'b0000000000;
    pxcRom[2797] <= 10'b0000000000;
    pxcRom[2798] <= 10'b0000000000;
    pxcRom[2799] <= 10'b0000000000;
    pxcRom[2800] <= 10'b0000000000;
    pxcRom[2801] <= 10'b0000000000;
    pxcRom[2802] <= 10'b0000000000;
    pxcRom[2803] <= 10'b0000000000;
    pxcRom[2804] <= 10'b0000000001;
    pxcRom[2805] <= 10'b0000000010;
    pxcRom[2806] <= 10'b0000000011;
    pxcRom[2807] <= 10'b0000000100;
    pxcRom[2808] <= 10'b0000000110;
    pxcRom[2809] <= 10'b0000001010;
    pxcRom[2810] <= 10'b0000001110;
    pxcRom[2811] <= 10'b0000010001;
    pxcRom[2812] <= 10'b0000010010;
    pxcRom[2813] <= 10'b0000010010;
    pxcRom[2814] <= 10'b0000010100;
    pxcRom[2815] <= 10'b0000011010;
    pxcRom[2816] <= 10'b0000101000;
    pxcRom[2817] <= 10'b0000111111;
    pxcRom[2818] <= 10'b0001001101;
    pxcRom[2819] <= 10'b0001000001;
    pxcRom[2820] <= 10'b0000101000;
    pxcRom[2821] <= 10'b0000010100;
    pxcRom[2822] <= 10'b0000001000;
    pxcRom[2823] <= 10'b0000000010;
    pxcRom[2824] <= 10'b0000000000;
    pxcRom[2825] <= 10'b0000000000;
    pxcRom[2826] <= 10'b0000000000;
    pxcRom[2827] <= 10'b0000000000;
    pxcRom[2828] <= 10'b0000000000;
    pxcRom[2829] <= 10'b0000000000;
    pxcRom[2830] <= 10'b0000000000;
    pxcRom[2831] <= 10'b0000000001;
    pxcRom[2832] <= 10'b0000000011;
    pxcRom[2833] <= 10'b0000000100;
    pxcRom[2834] <= 10'b0000000101;
    pxcRom[2835] <= 10'b0000000101;
    pxcRom[2836] <= 10'b0000000110;
    pxcRom[2837] <= 10'b0000000110;
    pxcRom[2838] <= 10'b0000000110;
    pxcRom[2839] <= 10'b0000000110;
    pxcRom[2840] <= 10'b0000000110;
    pxcRom[2841] <= 10'b0000000111;
    pxcRom[2842] <= 10'b0000001010;
    pxcRom[2843] <= 10'b0000010001;
    pxcRom[2844] <= 10'b0000100000;
    pxcRom[2845] <= 10'b0000110111;
    pxcRom[2846] <= 10'b0001001010;
    pxcRom[2847] <= 10'b0001000100;
    pxcRom[2848] <= 10'b0000101011;
    pxcRom[2849] <= 10'b0000010110;
    pxcRom[2850] <= 10'b0000001010;
    pxcRom[2851] <= 10'b0000000011;
    pxcRom[2852] <= 10'b0000000000;
    pxcRom[2853] <= 10'b0000000000;
    pxcRom[2854] <= 10'b0000000000;
    pxcRom[2855] <= 10'b0000000000;
    pxcRom[2856] <= 10'b0000000000;
    pxcRom[2857] <= 10'b0000000000;
    pxcRom[2858] <= 10'b0000000000;
    pxcRom[2859] <= 10'b0000000010;
    pxcRom[2860] <= 10'b0000000101;
    pxcRom[2861] <= 10'b0000001000;
    pxcRom[2862] <= 10'b0000001001;
    pxcRom[2863] <= 10'b0000001010;
    pxcRom[2864] <= 10'b0000001001;
    pxcRom[2865] <= 10'b0000001000;
    pxcRom[2866] <= 10'b0000000110;
    pxcRom[2867] <= 10'b0000000101;
    pxcRom[2868] <= 10'b0000000101;
    pxcRom[2869] <= 10'b0000000110;
    pxcRom[2870] <= 10'b0000001001;
    pxcRom[2871] <= 10'b0000010011;
    pxcRom[2872] <= 10'b0000100101;
    pxcRom[2873] <= 10'b0000111011;
    pxcRom[2874] <= 10'b0001001011;
    pxcRom[2875] <= 10'b0001000100;
    pxcRom[2876] <= 10'b0000101001;
    pxcRom[2877] <= 10'b0000010110;
    pxcRom[2878] <= 10'b0000001010;
    pxcRom[2879] <= 10'b0000000011;
    pxcRom[2880] <= 10'b0000000000;
    pxcRom[2881] <= 10'b0000000000;
    pxcRom[2882] <= 10'b0000000000;
    pxcRom[2883] <= 10'b0000000000;
    pxcRom[2884] <= 10'b0000000000;
    pxcRom[2885] <= 10'b0000000000;
    pxcRom[2886] <= 10'b0000000000;
    pxcRom[2887] <= 10'b0000000100;
    pxcRom[2888] <= 10'b0000001000;
    pxcRom[2889] <= 10'b0000001101;
    pxcRom[2890] <= 10'b0000010001;
    pxcRom[2891] <= 10'b0000010011;
    pxcRom[2892] <= 10'b0000010010;
    pxcRom[2893] <= 10'b0000010000;
    pxcRom[2894] <= 10'b0000001101;
    pxcRom[2895] <= 10'b0000001010;
    pxcRom[2896] <= 10'b0000001001;
    pxcRom[2897] <= 10'b0000001100;
    pxcRom[2898] <= 10'b0000010010;
    pxcRom[2899] <= 10'b0000011111;
    pxcRom[2900] <= 10'b0000110010;
    pxcRom[2901] <= 10'b0001001001;
    pxcRom[2902] <= 10'b0001001111;
    pxcRom[2903] <= 10'b0000111111;
    pxcRom[2904] <= 10'b0000100101;
    pxcRom[2905] <= 10'b0000010011;
    pxcRom[2906] <= 10'b0000001001;
    pxcRom[2907] <= 10'b0000000010;
    pxcRom[2908] <= 10'b0000000000;
    pxcRom[2909] <= 10'b0000000000;
    pxcRom[2910] <= 10'b0000000000;
    pxcRom[2911] <= 10'b0000000000;
    pxcRom[2912] <= 10'b0000000000;
    pxcRom[2913] <= 10'b0000000000;
    pxcRom[2914] <= 10'b0000000001;
    pxcRom[2915] <= 10'b0000000100;
    pxcRom[2916] <= 10'b0000001010;
    pxcRom[2917] <= 10'b0000010001;
    pxcRom[2918] <= 10'b0000011001;
    pxcRom[2919] <= 10'b0000011111;
    pxcRom[2920] <= 10'b0000100010;
    pxcRom[2921] <= 10'b0000100001;
    pxcRom[2922] <= 10'b0000011101;
    pxcRom[2923] <= 10'b0000011010;
    pxcRom[2924] <= 10'b0000011010;
    pxcRom[2925] <= 10'b0000011111;
    pxcRom[2926] <= 10'b0000101001;
    pxcRom[2927] <= 10'b0000111010;
    pxcRom[2928] <= 10'b0001001111;
    pxcRom[2929] <= 10'b0001011010;
    pxcRom[2930] <= 10'b0001001101;
    pxcRom[2931] <= 10'b0000110010;
    pxcRom[2932] <= 10'b0000011101;
    pxcRom[2933] <= 10'b0000001111;
    pxcRom[2934] <= 10'b0000000110;
    pxcRom[2935] <= 10'b0000000001;
    pxcRom[2936] <= 10'b0000000000;
    pxcRom[2937] <= 10'b0000000000;
    pxcRom[2938] <= 10'b0000000000;
    pxcRom[2939] <= 10'b0000000000;
    pxcRom[2940] <= 10'b0000000000;
    pxcRom[2941] <= 10'b0000000000;
    pxcRom[2942] <= 10'b0000000000;
    pxcRom[2943] <= 10'b0000000100;
    pxcRom[2944] <= 10'b0000001010;
    pxcRom[2945] <= 10'b0000010010;
    pxcRom[2946] <= 10'b0000011110;
    pxcRom[2947] <= 10'b0000101010;
    pxcRom[2948] <= 10'b0000110110;
    pxcRom[2949] <= 10'b0000111101;
    pxcRom[2950] <= 10'b0000111101;
    pxcRom[2951] <= 10'b0000111101;
    pxcRom[2952] <= 10'b0000111111;
    pxcRom[2953] <= 10'b0001000111;
    pxcRom[2954] <= 10'b0001010100;
    pxcRom[2955] <= 10'b0001100011;
    pxcRom[2956] <= 10'b0001101000;
    pxcRom[2957] <= 10'b0001010110;
    pxcRom[2958] <= 10'b0000111010;
    pxcRom[2959] <= 10'b0000100011;
    pxcRom[2960] <= 10'b0000010011;
    pxcRom[2961] <= 10'b0000001001;
    pxcRom[2962] <= 10'b0000000011;
    pxcRom[2963] <= 10'b0000000000;
    pxcRom[2964] <= 10'b0000000000;
    pxcRom[2965] <= 10'b0000000000;
    pxcRom[2966] <= 10'b0000000000;
    pxcRom[2967] <= 10'b0000000000;
    pxcRom[2968] <= 10'b0000000000;
    pxcRom[2969] <= 10'b0000000000;
    pxcRom[2970] <= 10'b0000000000;
    pxcRom[2971] <= 10'b0000000011;
    pxcRom[2972] <= 10'b0000000111;
    pxcRom[2973] <= 10'b0000001110;
    pxcRom[2974] <= 10'b0000011011;
    pxcRom[2975] <= 10'b0000101010;
    pxcRom[2976] <= 10'b0000111110;
    pxcRom[2977] <= 10'b0001010010;
    pxcRom[2978] <= 10'b0001100010;
    pxcRom[2979] <= 10'b0001101101;
    pxcRom[2980] <= 10'b0001110100;
    pxcRom[2981] <= 10'b0001111010;
    pxcRom[2982] <= 10'b0001111001;
    pxcRom[2983] <= 10'b0001101101;
    pxcRom[2984] <= 10'b0001010101;
    pxcRom[2985] <= 10'b0000111001;
    pxcRom[2986] <= 10'b0000100011;
    pxcRom[2987] <= 10'b0000010011;
    pxcRom[2988] <= 10'b0000001001;
    pxcRom[2989] <= 10'b0000000100;
    pxcRom[2990] <= 10'b0000000001;
    pxcRom[2991] <= 10'b0000000000;
    pxcRom[2992] <= 10'b0000000000;
    pxcRom[2993] <= 10'b0000000000;
    pxcRom[2994] <= 10'b0000000000;
    pxcRom[2995] <= 10'b0000000000;
    pxcRom[2996] <= 10'b0000000000;
    pxcRom[2997] <= 10'b0000000000;
    pxcRom[2998] <= 10'b0000000000;
    pxcRom[2999] <= 10'b0000000001;
    pxcRom[3000] <= 10'b0000000100;
    pxcRom[3001] <= 10'b0000001000;
    pxcRom[3002] <= 10'b0000010000;
    pxcRom[3003] <= 10'b0000011100;
    pxcRom[3004] <= 10'b0000101100;
    pxcRom[3005] <= 10'b0000111110;
    pxcRom[3006] <= 10'b0001010001;
    pxcRom[3007] <= 10'b0001100000;
    pxcRom[3008] <= 10'b0001100111;
    pxcRom[3009] <= 10'b0001100001;
    pxcRom[3010] <= 10'b0001010010;
    pxcRom[3011] <= 10'b0000111111;
    pxcRom[3012] <= 10'b0000101011;
    pxcRom[3013] <= 10'b0000011011;
    pxcRom[3014] <= 10'b0000001111;
    pxcRom[3015] <= 10'b0000001000;
    pxcRom[3016] <= 10'b0000000011;
    pxcRom[3017] <= 10'b0000000001;
    pxcRom[3018] <= 10'b0000000000;
    pxcRom[3019] <= 10'b0000000000;
    pxcRom[3020] <= 10'b0000000000;
    pxcRom[3021] <= 10'b0000000000;
    pxcRom[3022] <= 10'b0000000000;
    pxcRom[3023] <= 10'b0000000000;
    pxcRom[3024] <= 10'b0000000000;
    pxcRom[3025] <= 10'b0000000000;
    pxcRom[3026] <= 10'b0000000000;
    pxcRom[3027] <= 10'b0000000000;
    pxcRom[3028] <= 10'b0000000001;
    pxcRom[3029] <= 10'b0000000011;
    pxcRom[3030] <= 10'b0000000110;
    pxcRom[3031] <= 10'b0000001010;
    pxcRom[3032] <= 10'b0000001111;
    pxcRom[3033] <= 10'b0000010101;
    pxcRom[3034] <= 10'b0000011011;
    pxcRom[3035] <= 10'b0000011111;
    pxcRom[3036] <= 10'b0000100000;
    pxcRom[3037] <= 10'b0000011110;
    pxcRom[3038] <= 10'b0000011001;
    pxcRom[3039] <= 10'b0000010011;
    pxcRom[3040] <= 10'b0000001100;
    pxcRom[3041] <= 10'b0000000111;
    pxcRom[3042] <= 10'b0000000100;
    pxcRom[3043] <= 10'b0000000001;
    pxcRom[3044] <= 10'b0000000000;
    pxcRom[3045] <= 10'b0000000000;
    pxcRom[3046] <= 10'b0000000000;
    pxcRom[3047] <= 10'b0000000000;
    pxcRom[3048] <= 10'b0000000000;
    pxcRom[3049] <= 10'b0000000000;
    pxcRom[3050] <= 10'b0000000000;
    pxcRom[3051] <= 10'b0000000000;
    pxcRom[3052] <= 10'b0000000000;
    pxcRom[3053] <= 10'b0000000000;
    pxcRom[3054] <= 10'b0000000000;
    pxcRom[3055] <= 10'b0000000000;
    pxcRom[3056] <= 10'b0000000000;
    pxcRom[3057] <= 10'b0000000000;
    pxcRom[3058] <= 10'b0000000000;
    pxcRom[3059] <= 10'b0000000001;
    pxcRom[3060] <= 10'b0000000001;
    pxcRom[3061] <= 10'b0000000010;
    pxcRom[3062] <= 10'b0000000010;
    pxcRom[3063] <= 10'b0000000011;
    pxcRom[3064] <= 10'b0000000011;
    pxcRom[3065] <= 10'b0000000011;
    pxcRom[3066] <= 10'b0000000010;
    pxcRom[3067] <= 10'b0000000010;
    pxcRom[3068] <= 10'b0000000001;
    pxcRom[3069] <= 10'b0000000000;
    pxcRom[3070] <= 10'b0000000000;
    pxcRom[3071] <= 10'b0000000000;
    pxcRom[3072] <= 10'b0000000000;
    pxcRom[3073] <= 10'b0000000000;
    pxcRom[3074] <= 10'b0000000000;
    pxcRom[3075] <= 10'b0000000000;
    pxcRom[3076] <= 10'b0000000000;
    pxcRom[3077] <= 10'b0000000000;
    pxcRom[3078] <= 10'b0000000000;
    pxcRom[3079] <= 10'b0000000000;
    pxcRom[3080] <= 10'b0000000000;
    pxcRom[3081] <= 10'b0000000000;
    pxcRom[3082] <= 10'b0000000000;
    pxcRom[3083] <= 10'b0000000000;
    pxcRom[3084] <= 10'b0000000000;
    pxcRom[3085] <= 10'b0000000000;
    pxcRom[3086] <= 10'b0000000000;
    pxcRom[3087] <= 10'b0000000000;
    pxcRom[3088] <= 10'b0000000000;
    pxcRom[3089] <= 10'b0000000000;
    pxcRom[3090] <= 10'b0000000000;
    pxcRom[3091] <= 10'b0000000000;
    pxcRom[3092] <= 10'b0000000000;
    pxcRom[3093] <= 10'b0000000000;
    pxcRom[3094] <= 10'b0000000000;
    pxcRom[3095] <= 10'b0000000000;
    pxcRom[3096] <= 10'b0000000000;
    pxcRom[3097] <= 10'b0000000000;
    pxcRom[3098] <= 10'b0000000000;
    pxcRom[3099] <= 10'b0000000000;
    pxcRom[3100] <= 10'b0000000000;
    pxcRom[3101] <= 10'b0000000000;
    pxcRom[3102] <= 10'b0000000000;
    pxcRom[3103] <= 10'b0000000000;
    pxcRom[3104] <= 10'b0000000000;
    pxcRom[3105] <= 10'b0000000000;
    pxcRom[3106] <= 10'b0000000000;
    pxcRom[3107] <= 10'b0000000000;
    pxcRom[3108] <= 10'b0000000000;
    pxcRom[3109] <= 10'b0000000000;
    pxcRom[3110] <= 10'b0000000000;
    pxcRom[3111] <= 10'b0000000000;
    pxcRom[3112] <= 10'b0000000000;
    pxcRom[3113] <= 10'b0000000000;
    pxcRom[3114] <= 10'b0000000000;
    pxcRom[3115] <= 10'b0000000000;
    pxcRom[3116] <= 10'b0000000000;
    pxcRom[3117] <= 10'b0000000000;
    pxcRom[3118] <= 10'b0000000000;
    pxcRom[3119] <= 10'b0000000000;
    pxcRom[3120] <= 10'b0000000000;
    pxcRom[3121] <= 10'b0000000000;
    pxcRom[3122] <= 10'b0000000000;
    pxcRom[3123] <= 10'b0000000000;
    pxcRom[3124] <= 10'b0000000000;
    pxcRom[3125] <= 10'b0000000000;
    pxcRom[3126] <= 10'b0000000000;
    pxcRom[3127] <= 10'b0000000000;
    pxcRom[3128] <= 10'b0000000000;
    pxcRom[3129] <= 10'b0000000000;
    pxcRom[3130] <= 10'b0000000000;
    pxcRom[3131] <= 10'b0000000000;
    pxcRom[3132] <= 10'b0000000000;
    pxcRom[3133] <= 10'b0000000000;
    pxcRom[3134] <= 10'b0000000000;
    pxcRom[3135] <= 10'b0000000000;
    pxcRom[3136] <= 10'b0000000000;
    pxcRom[3137] <= 10'b0000000000;
    pxcRom[3138] <= 10'b0000000000;
    pxcRom[3139] <= 10'b0000000000;
    pxcRom[3140] <= 10'b0000000000;
    pxcRom[3141] <= 10'b0000000000;
    pxcRom[3142] <= 10'b0000000000;
    pxcRom[3143] <= 10'b0000000000;
    pxcRom[3144] <= 10'b0000000000;
    pxcRom[3145] <= 10'b0000000000;
    pxcRom[3146] <= 10'b0000000000;
    pxcRom[3147] <= 10'b0000000000;
    pxcRom[3148] <= 10'b0000000000;
    pxcRom[3149] <= 10'b0000000000;
    pxcRom[3150] <= 10'b0000000000;
    pxcRom[3151] <= 10'b0000000000;
    pxcRom[3152] <= 10'b0000000000;
    pxcRom[3153] <= 10'b0000000000;
    pxcRom[3154] <= 10'b0000000000;
    pxcRom[3155] <= 10'b0000000000;
    pxcRom[3156] <= 10'b0000000000;
    pxcRom[3157] <= 10'b0000000000;
    pxcRom[3158] <= 10'b0000000000;
    pxcRom[3159] <= 10'b0000000000;
    pxcRom[3160] <= 10'b0000000000;
    pxcRom[3161] <= 10'b0000000000;
    pxcRom[3162] <= 10'b0000000000;
    pxcRom[3163] <= 10'b0000000000;
    pxcRom[3164] <= 10'b0000000000;
    pxcRom[3165] <= 10'b0000000000;
    pxcRom[3166] <= 10'b0000000000;
    pxcRom[3167] <= 10'b0000000000;
    pxcRom[3168] <= 10'b0000000000;
    pxcRom[3169] <= 10'b0000000000;
    pxcRom[3170] <= 10'b0000000000;
    pxcRom[3171] <= 10'b0000000000;
    pxcRom[3172] <= 10'b0000000000;
    pxcRom[3173] <= 10'b0000000000;
    pxcRom[3174] <= 10'b0000000000;
    pxcRom[3175] <= 10'b0000000000;
    pxcRom[3176] <= 10'b0000000000;
    pxcRom[3177] <= 10'b0000000000;
    pxcRom[3178] <= 10'b0000000000;
    pxcRom[3179] <= 10'b0000000000;
    pxcRom[3180] <= 10'b0000000000;
    pxcRom[3181] <= 10'b0000000000;
    pxcRom[3182] <= 10'b0000000000;
    pxcRom[3183] <= 10'b0000000000;
    pxcRom[3184] <= 10'b0000000000;
    pxcRom[3185] <= 10'b0000000000;
    pxcRom[3186] <= 10'b0000000000;
    pxcRom[3187] <= 10'b0000000000;
    pxcRom[3188] <= 10'b0000000000;
    pxcRom[3189] <= 10'b0000000000;
    pxcRom[3190] <= 10'b0000000000;
    pxcRom[3191] <= 10'b0000000000;
    pxcRom[3192] <= 10'b0000000000;
    pxcRom[3193] <= 10'b0000000000;
    pxcRom[3194] <= 10'b0000000000;
    pxcRom[3195] <= 10'b0000000000;
    pxcRom[3196] <= 10'b0000000000;
    pxcRom[3197] <= 10'b0000000000;
    pxcRom[3198] <= 10'b0000000000;
    pxcRom[3199] <= 10'b0000000000;
    pxcRom[3200] <= 10'b0000000000;
    pxcRom[3201] <= 10'b0000000000;
    pxcRom[3202] <= 10'b0000000000;
    pxcRom[3203] <= 10'b0000000000;
    pxcRom[3204] <= 10'b0000000000;
    pxcRom[3205] <= 10'b0000000000;
    pxcRom[3206] <= 10'b0000000000;
    pxcRom[3207] <= 10'b0000000000;
    pxcRom[3208] <= 10'b0000000000;
    pxcRom[3209] <= 10'b0000000000;
    pxcRom[3210] <= 10'b0000000000;
    pxcRom[3211] <= 10'b0000000000;
    pxcRom[3212] <= 10'b0000000000;
    pxcRom[3213] <= 10'b0000000000;
    pxcRom[3214] <= 10'b0000000000;
    pxcRom[3215] <= 10'b0000000000;
    pxcRom[3216] <= 10'b0000000000;
    pxcRom[3217] <= 10'b0000000000;
    pxcRom[3218] <= 10'b0000000000;
    pxcRom[3219] <= 10'b0000000000;
    pxcRom[3220] <= 10'b0000000000;
    pxcRom[3221] <= 10'b0000000000;
    pxcRom[3222] <= 10'b0000000000;
    pxcRom[3223] <= 10'b0000000000;
    pxcRom[3224] <= 10'b0000000000;
    pxcRom[3225] <= 10'b0000000000;
    pxcRom[3226] <= 10'b0000000000;
    pxcRom[3227] <= 10'b0000000000;
    pxcRom[3228] <= 10'b0000000000;
    pxcRom[3229] <= 10'b0000000000;
    pxcRom[3230] <= 10'b0000000000;
    pxcRom[3231] <= 10'b0000000000;
    pxcRom[3232] <= 10'b0000000000;
    pxcRom[3233] <= 10'b0000000000;
    pxcRom[3234] <= 10'b0000000000;
    pxcRom[3235] <= 10'b0000000000;
    pxcRom[3236] <= 10'b0000000000;
    pxcRom[3237] <= 10'b0000000000;
    pxcRom[3238] <= 10'b0000000000;
    pxcRom[3239] <= 10'b0000000000;
    pxcRom[3240] <= 10'b0000000000;
    pxcRom[3241] <= 10'b0000000000;
    pxcRom[3242] <= 10'b0000000000;
    pxcRom[3243] <= 10'b0000000000;
    pxcRom[3244] <= 10'b0000000000;
    pxcRom[3245] <= 10'b0000000000;
    pxcRom[3246] <= 10'b0000000000;
    pxcRom[3247] <= 10'b0000000000;
    pxcRom[3248] <= 10'b0000000000;
    pxcRom[3249] <= 10'b0000000000;
    pxcRom[3250] <= 10'b0000000000;
    pxcRom[3251] <= 10'b0000000000;
    pxcRom[3252] <= 10'b0000000000;
    pxcRom[3253] <= 10'b0000000000;
    pxcRom[3254] <= 10'b0000000000;
    pxcRom[3255] <= 10'b0000000000;
    pxcRom[3256] <= 10'b0000000000;
    pxcRom[3257] <= 10'b0000000000;
    pxcRom[3258] <= 10'b0000000001;
    pxcRom[3259] <= 10'b0000000001;
    pxcRom[3260] <= 10'b0000000001;
    pxcRom[3261] <= 10'b0000000001;
    pxcRom[3262] <= 10'b0000000001;
    pxcRom[3263] <= 10'b0000000001;
    pxcRom[3264] <= 10'b0000000010;
    pxcRom[3265] <= 10'b0000000011;
    pxcRom[3266] <= 10'b0000000011;
    pxcRom[3267] <= 10'b0000000100;
    pxcRom[3268] <= 10'b0000000100;
    pxcRom[3269] <= 10'b0000000100;
    pxcRom[3270] <= 10'b0000000011;
    pxcRom[3271] <= 10'b0000000001;
    pxcRom[3272] <= 10'b0000000000;
    pxcRom[3273] <= 10'b0000000000;
    pxcRom[3274] <= 10'b0000000000;
    pxcRom[3275] <= 10'b0000000000;
    pxcRom[3276] <= 10'b0000000000;
    pxcRom[3277] <= 10'b0000000000;
    pxcRom[3278] <= 10'b0000000000;
    pxcRom[3279] <= 10'b0000000000;
    pxcRom[3280] <= 10'b0000000000;
    pxcRom[3281] <= 10'b0000000000;
    pxcRom[3282] <= 10'b0000000001;
    pxcRom[3283] <= 10'b0000000010;
    pxcRom[3284] <= 10'b0000000011;
    pxcRom[3285] <= 10'b0000000101;
    pxcRom[3286] <= 10'b0000000111;
    pxcRom[3287] <= 10'b0000000111;
    pxcRom[3288] <= 10'b0000001000;
    pxcRom[3289] <= 10'b0000000111;
    pxcRom[3290] <= 10'b0000000110;
    pxcRom[3291] <= 10'b0000000110;
    pxcRom[3292] <= 10'b0000001001;
    pxcRom[3293] <= 10'b0000001100;
    pxcRom[3294] <= 10'b0000010000;
    pxcRom[3295] <= 10'b0000010001;
    pxcRom[3296] <= 10'b0000010000;
    pxcRom[3297] <= 10'b0000001101;
    pxcRom[3298] <= 10'b0000001010;
    pxcRom[3299] <= 10'b0000000110;
    pxcRom[3300] <= 10'b0000000011;
    pxcRom[3301] <= 10'b0000000000;
    pxcRom[3302] <= 10'b0000000000;
    pxcRom[3303] <= 10'b0000000000;
    pxcRom[3304] <= 10'b0000000000;
    pxcRom[3305] <= 10'b0000000000;
    pxcRom[3306] <= 10'b0000000000;
    pxcRom[3307] <= 10'b0000000000;
    pxcRom[3308] <= 10'b0000000000;
    pxcRom[3309] <= 10'b0000000001;
    pxcRom[3310] <= 10'b0000000010;
    pxcRom[3311] <= 10'b0000000100;
    pxcRom[3312] <= 10'b0000001000;
    pxcRom[3313] <= 10'b0000001100;
    pxcRom[3314] <= 10'b0000010000;
    pxcRom[3315] <= 10'b0000010010;
    pxcRom[3316] <= 10'b0000010001;
    pxcRom[3317] <= 10'b0000001110;
    pxcRom[3318] <= 10'b0000001011;
    pxcRom[3319] <= 10'b0000001011;
    pxcRom[3320] <= 10'b0000001111;
    pxcRom[3321] <= 10'b0000010110;
    pxcRom[3322] <= 10'b0000011101;
    pxcRom[3323] <= 10'b0000011110;
    pxcRom[3324] <= 10'b0000011011;
    pxcRom[3325] <= 10'b0000010101;
    pxcRom[3326] <= 10'b0000001111;
    pxcRom[3327] <= 10'b0000001001;
    pxcRom[3328] <= 10'b0000000100;
    pxcRom[3329] <= 10'b0000000001;
    pxcRom[3330] <= 10'b0000000000;
    pxcRom[3331] <= 10'b0000000000;
    pxcRom[3332] <= 10'b0000000000;
    pxcRom[3333] <= 10'b0000000000;
    pxcRom[3334] <= 10'b0000000000;
    pxcRom[3335] <= 10'b0000000000;
    pxcRom[3336] <= 10'b0000000000;
    pxcRom[3337] <= 10'b0000000010;
    pxcRom[3338] <= 10'b0000000100;
    pxcRom[3339] <= 10'b0000000111;
    pxcRom[3340] <= 10'b0000001101;
    pxcRom[3341] <= 10'b0000010101;
    pxcRom[3342] <= 10'b0000011011;
    pxcRom[3343] <= 10'b0000011101;
    pxcRom[3344] <= 10'b0000011010;
    pxcRom[3345] <= 10'b0000010101;
    pxcRom[3346] <= 10'b0000001111;
    pxcRom[3347] <= 10'b0000001101;
    pxcRom[3348] <= 10'b0000010011;
    pxcRom[3349] <= 10'b0000011110;
    pxcRom[3350] <= 10'b0000101000;
    pxcRom[3351] <= 10'b0000101010;
    pxcRom[3352] <= 10'b0000100011;
    pxcRom[3353] <= 10'b0000011001;
    pxcRom[3354] <= 10'b0000010000;
    pxcRom[3355] <= 10'b0000001001;
    pxcRom[3356] <= 10'b0000000100;
    pxcRom[3357] <= 10'b0000000001;
    pxcRom[3358] <= 10'b0000000000;
    pxcRom[3359] <= 10'b0000000000;
    pxcRom[3360] <= 10'b0000000000;
    pxcRom[3361] <= 10'b0000000000;
    pxcRom[3362] <= 10'b0000000000;
    pxcRom[3363] <= 10'b0000000000;
    pxcRom[3364] <= 10'b0000000001;
    pxcRom[3365] <= 10'b0000000010;
    pxcRom[3366] <= 10'b0000000101;
    pxcRom[3367] <= 10'b0000001010;
    pxcRom[3368] <= 10'b0000010011;
    pxcRom[3369] <= 10'b0000011110;
    pxcRom[3370] <= 10'b0000100111;
    pxcRom[3371] <= 10'b0000101001;
    pxcRom[3372] <= 10'b0000100100;
    pxcRom[3373] <= 10'b0000011001;
    pxcRom[3374] <= 10'b0000010000;
    pxcRom[3375] <= 10'b0000001110;
    pxcRom[3376] <= 10'b0000010110;
    pxcRom[3377] <= 10'b0000100110;
    pxcRom[3378] <= 10'b0000110101;
    pxcRom[3379] <= 10'b0000110101;
    pxcRom[3380] <= 10'b0000101000;
    pxcRom[3381] <= 10'b0000011001;
    pxcRom[3382] <= 10'b0000001110;
    pxcRom[3383] <= 10'b0000000111;
    pxcRom[3384] <= 10'b0000000010;
    pxcRom[3385] <= 10'b0000000000;
    pxcRom[3386] <= 10'b0000000000;
    pxcRom[3387] <= 10'b0000000000;
    pxcRom[3388] <= 10'b0000000000;
    pxcRom[3389] <= 10'b0000000000;
    pxcRom[3390] <= 10'b0000000000;
    pxcRom[3391] <= 10'b0000000000;
    pxcRom[3392] <= 10'b0000000001;
    pxcRom[3393] <= 10'b0000000010;
    pxcRom[3394] <= 10'b0000000110;
    pxcRom[3395] <= 10'b0000001110;
    pxcRom[3396] <= 10'b0000011001;
    pxcRom[3397] <= 10'b0000101001;
    pxcRom[3398] <= 10'b0000110100;
    pxcRom[3399] <= 10'b0000110100;
    pxcRom[3400] <= 10'b0000100111;
    pxcRom[3401] <= 10'b0000011001;
    pxcRom[3402] <= 10'b0000001110;
    pxcRom[3403] <= 10'b0000001110;
    pxcRom[3404] <= 10'b0000011001;
    pxcRom[3405] <= 10'b0000110000;
    pxcRom[3406] <= 10'b0001000010;
    pxcRom[3407] <= 10'b0000111110;
    pxcRom[3408] <= 10'b0000101001;
    pxcRom[3409] <= 10'b0000010110;
    pxcRom[3410] <= 10'b0000001100;
    pxcRom[3411] <= 10'b0000000100;
    pxcRom[3412] <= 10'b0000000001;
    pxcRom[3413] <= 10'b0000000000;
    pxcRom[3414] <= 10'b0000000000;
    pxcRom[3415] <= 10'b0000000000;
    pxcRom[3416] <= 10'b0000000000;
    pxcRom[3417] <= 10'b0000000000;
    pxcRom[3418] <= 10'b0000000000;
    pxcRom[3419] <= 10'b0000000000;
    pxcRom[3420] <= 10'b0000000001;
    pxcRom[3421] <= 10'b0000000011;
    pxcRom[3422] <= 10'b0000001000;
    pxcRom[3423] <= 10'b0000010010;
    pxcRom[3424] <= 10'b0000100011;
    pxcRom[3425] <= 10'b0000110111;
    pxcRom[3426] <= 10'b0001000010;
    pxcRom[3427] <= 10'b0000111000;
    pxcRom[3428] <= 10'b0000100101;
    pxcRom[3429] <= 10'b0000010100;
    pxcRom[3430] <= 10'b0000001010;
    pxcRom[3431] <= 10'b0000001101;
    pxcRom[3432] <= 10'b0000100000;
    pxcRom[3433] <= 10'b0000111110;
    pxcRom[3434] <= 10'b0001010010;
    pxcRom[3435] <= 10'b0001000000;
    pxcRom[3436] <= 10'b0000100101;
    pxcRom[3437] <= 10'b0000010010;
    pxcRom[3438] <= 10'b0000001000;
    pxcRom[3439] <= 10'b0000000010;
    pxcRom[3440] <= 10'b0000000000;
    pxcRom[3441] <= 10'b0000000000;
    pxcRom[3442] <= 10'b0000000000;
    pxcRom[3443] <= 10'b0000000000;
    pxcRom[3444] <= 10'b0000000000;
    pxcRom[3445] <= 10'b0000000000;
    pxcRom[3446] <= 10'b0000000000;
    pxcRom[3447] <= 10'b0000000000;
    pxcRom[3448] <= 10'b0000000001;
    pxcRom[3449] <= 10'b0000000100;
    pxcRom[3450] <= 10'b0000001100;
    pxcRom[3451] <= 10'b0000011010;
    pxcRom[3452] <= 10'b0000110000;
    pxcRom[3453] <= 10'b0001001001;
    pxcRom[3454] <= 10'b0001001100;
    pxcRom[3455] <= 10'b0000110101;
    pxcRom[3456] <= 10'b0000011101;
    pxcRom[3457] <= 10'b0000001101;
    pxcRom[3458] <= 10'b0000000111;
    pxcRom[3459] <= 10'b0000010000;
    pxcRom[3460] <= 10'b0000101011;
    pxcRom[3461] <= 10'b0001010010;
    pxcRom[3462] <= 10'b0001011110;
    pxcRom[3463] <= 10'b0000111101;
    pxcRom[3464] <= 10'b0000011111;
    pxcRom[3465] <= 10'b0000001101;
    pxcRom[3466] <= 10'b0000000101;
    pxcRom[3467] <= 10'b0000000001;
    pxcRom[3468] <= 10'b0000000000;
    pxcRom[3469] <= 10'b0000000000;
    pxcRom[3470] <= 10'b0000000000;
    pxcRom[3471] <= 10'b0000000000;
    pxcRom[3472] <= 10'b0000000000;
    pxcRom[3473] <= 10'b0000000000;
    pxcRom[3474] <= 10'b0000000000;
    pxcRom[3475] <= 10'b0000000000;
    pxcRom[3476] <= 10'b0000000001;
    pxcRom[3477] <= 10'b0000000110;
    pxcRom[3478] <= 10'b0000010000;
    pxcRom[3479] <= 10'b0000100100;
    pxcRom[3480] <= 10'b0001000010;
    pxcRom[3481] <= 10'b0001011100;
    pxcRom[3482] <= 10'b0001010000;
    pxcRom[3483] <= 10'b0000110000;
    pxcRom[3484] <= 10'b0000011000;
    pxcRom[3485] <= 10'b0000001100;
    pxcRom[3486] <= 10'b0000001011;
    pxcRom[3487] <= 10'b0000011010;
    pxcRom[3488] <= 10'b0000111111;
    pxcRom[3489] <= 10'b0001101100;
    pxcRom[3490] <= 10'b0001100010;
    pxcRom[3491] <= 10'b0000111001;
    pxcRom[3492] <= 10'b0000011011;
    pxcRom[3493] <= 10'b0000001100;
    pxcRom[3494] <= 10'b0000000101;
    pxcRom[3495] <= 10'b0000000001;
    pxcRom[3496] <= 10'b0000000000;
    pxcRom[3497] <= 10'b0000000000;
    pxcRom[3498] <= 10'b0000000000;
    pxcRom[3499] <= 10'b0000000000;
    pxcRom[3500] <= 10'b0000000000;
    pxcRom[3501] <= 10'b0000000000;
    pxcRom[3502] <= 10'b0000000000;
    pxcRom[3503] <= 10'b0000000000;
    pxcRom[3504] <= 10'b0000000010;
    pxcRom[3505] <= 10'b0000001000;
    pxcRom[3506] <= 10'b0000010111;
    pxcRom[3507] <= 10'b0000110000;
    pxcRom[3508] <= 10'b0001010110;
    pxcRom[3509] <= 10'b0001101111;
    pxcRom[3510] <= 10'b0001010101;
    pxcRom[3511] <= 10'b0000110010;
    pxcRom[3512] <= 10'b0000011101;
    pxcRom[3513] <= 10'b0000010110;
    pxcRom[3514] <= 10'b0000011010;
    pxcRom[3515] <= 10'b0000110001;
    pxcRom[3516] <= 10'b0001011110;
    pxcRom[3517] <= 10'b0010000111;
    pxcRom[3518] <= 10'b0001100100;
    pxcRom[3519] <= 10'b0000111000;
    pxcRom[3520] <= 10'b0000011100;
    pxcRom[3521] <= 10'b0000001110;
    pxcRom[3522] <= 10'b0000000110;
    pxcRom[3523] <= 10'b0000000011;
    pxcRom[3524] <= 10'b0000000001;
    pxcRom[3525] <= 10'b0000000000;
    pxcRom[3526] <= 10'b0000000000;
    pxcRom[3527] <= 10'b0000000000;
    pxcRom[3528] <= 10'b0000000000;
    pxcRom[3529] <= 10'b0000000000;
    pxcRom[3530] <= 10'b0000000000;
    pxcRom[3531] <= 10'b0000000000;
    pxcRom[3532] <= 10'b0000000011;
    pxcRom[3533] <= 10'b0000001011;
    pxcRom[3534] <= 10'b0000011110;
    pxcRom[3535] <= 10'b0000111100;
    pxcRom[3536] <= 10'b0001100110;
    pxcRom[3537] <= 10'b0001111011;
    pxcRom[3538] <= 10'b0001100110;
    pxcRom[3539] <= 10'b0001000110;
    pxcRom[3540] <= 10'b0000111000;
    pxcRom[3541] <= 10'b0000110101;
    pxcRom[3542] <= 10'b0000111110;
    pxcRom[3543] <= 10'b0001011010;
    pxcRom[3544] <= 10'b0010001011;
    pxcRom[3545] <= 10'b0010011101;
    pxcRom[3546] <= 10'b0001101010;
    pxcRom[3547] <= 10'b0000111011;
    pxcRom[3548] <= 10'b0000100000;
    pxcRom[3549] <= 10'b0000010001;
    pxcRom[3550] <= 10'b0000001001;
    pxcRom[3551] <= 10'b0000000100;
    pxcRom[3552] <= 10'b0000000001;
    pxcRom[3553] <= 10'b0000000000;
    pxcRom[3554] <= 10'b0000000000;
    pxcRom[3555] <= 10'b0000000000;
    pxcRom[3556] <= 10'b0000000000;
    pxcRom[3557] <= 10'b0000000000;
    pxcRom[3558] <= 10'b0000000000;
    pxcRom[3559] <= 10'b0000000000;
    pxcRom[3560] <= 10'b0000000011;
    pxcRom[3561] <= 10'b0000001101;
    pxcRom[3562] <= 10'b0000100000;
    pxcRom[3563] <= 10'b0000111101;
    pxcRom[3564] <= 10'b0001100001;
    pxcRom[3565] <= 10'b0001111011;
    pxcRom[3566] <= 10'b0001110111;
    pxcRom[3567] <= 10'b0001100111;
    pxcRom[3568] <= 10'b0001100000;
    pxcRom[3569] <= 10'b0001100001;
    pxcRom[3570] <= 10'b0001110000;
    pxcRom[3571] <= 10'b0010001011;
    pxcRom[3572] <= 10'b0010110011;
    pxcRom[3573] <= 10'b0010100110;
    pxcRom[3574] <= 10'b0001101000;
    pxcRom[3575] <= 10'b0000111011;
    pxcRom[3576] <= 10'b0000100000;
    pxcRom[3577] <= 10'b0000010001;
    pxcRom[3578] <= 10'b0000001001;
    pxcRom[3579] <= 10'b0000000101;
    pxcRom[3580] <= 10'b0000000010;
    pxcRom[3581] <= 10'b0000000000;
    pxcRom[3582] <= 10'b0000000000;
    pxcRom[3583] <= 10'b0000000000;
    pxcRom[3584] <= 10'b0000000000;
    pxcRom[3585] <= 10'b0000000000;
    pxcRom[3586] <= 10'b0000000000;
    pxcRom[3587] <= 10'b0000000000;
    pxcRom[3588] <= 10'b0000000011;
    pxcRom[3589] <= 10'b0000001101;
    pxcRom[3590] <= 10'b0000011100;
    pxcRom[3591] <= 10'b0000101111;
    pxcRom[3592] <= 10'b0001000110;
    pxcRom[3593] <= 10'b0001010110;
    pxcRom[3594] <= 10'b0001011100;
    pxcRom[3595] <= 10'b0001011101;
    pxcRom[3596] <= 10'b0001011110;
    pxcRom[3597] <= 10'b0001100100;
    pxcRom[3598] <= 10'b0001110100;
    pxcRom[3599] <= 10'b0010010000;
    pxcRom[3600] <= 10'b0010100111;
    pxcRom[3601] <= 10'b0010000011;
    pxcRom[3602] <= 10'b0001010000;
    pxcRom[3603] <= 10'b0000101101;
    pxcRom[3604] <= 10'b0000011000;
    pxcRom[3605] <= 10'b0000001101;
    pxcRom[3606] <= 10'b0000000111;
    pxcRom[3607] <= 10'b0000000011;
    pxcRom[3608] <= 10'b0000000001;
    pxcRom[3609] <= 10'b0000000000;
    pxcRom[3610] <= 10'b0000000000;
    pxcRom[3611] <= 10'b0000000000;
    pxcRom[3612] <= 10'b0000000000;
    pxcRom[3613] <= 10'b0000000000;
    pxcRom[3614] <= 10'b0000000000;
    pxcRom[3615] <= 10'b0000000000;
    pxcRom[3616] <= 10'b0000000010;
    pxcRom[3617] <= 10'b0000001000;
    pxcRom[3618] <= 10'b0000010010;
    pxcRom[3619] <= 10'b0000011100;
    pxcRom[3620] <= 10'b0000100101;
    pxcRom[3621] <= 10'b0000101011;
    pxcRom[3622] <= 10'b0000101101;
    pxcRom[3623] <= 10'b0000110001;
    pxcRom[3624] <= 10'b0000110101;
    pxcRom[3625] <= 10'b0000111111;
    pxcRom[3626] <= 10'b0001010011;
    pxcRom[3627] <= 10'b0001101100;
    pxcRom[3628] <= 10'b0001110101;
    pxcRom[3629] <= 10'b0001010101;
    pxcRom[3630] <= 10'b0000110011;
    pxcRom[3631] <= 10'b0000011100;
    pxcRom[3632] <= 10'b0000001111;
    pxcRom[3633] <= 10'b0000001000;
    pxcRom[3634] <= 10'b0000000100;
    pxcRom[3635] <= 10'b0000000010;
    pxcRom[3636] <= 10'b0000000000;
    pxcRom[3637] <= 10'b0000000000;
    pxcRom[3638] <= 10'b0000000000;
    pxcRom[3639] <= 10'b0000000000;
    pxcRom[3640] <= 10'b0000000000;
    pxcRom[3641] <= 10'b0000000000;
    pxcRom[3642] <= 10'b0000000000;
    pxcRom[3643] <= 10'b0000000000;
    pxcRom[3644] <= 10'b0000000001;
    pxcRom[3645] <= 10'b0000000100;
    pxcRom[3646] <= 10'b0000001000;
    pxcRom[3647] <= 10'b0000001100;
    pxcRom[3648] <= 10'b0000001111;
    pxcRom[3649] <= 10'b0000010001;
    pxcRom[3650] <= 10'b0000010010;
    pxcRom[3651] <= 10'b0000010101;
    pxcRom[3652] <= 10'b0000011100;
    pxcRom[3653] <= 10'b0000101001;
    pxcRom[3654] <= 10'b0000111100;
    pxcRom[3655] <= 10'b0001001110;
    pxcRom[3656] <= 10'b0001001101;
    pxcRom[3657] <= 10'b0000110111;
    pxcRom[3658] <= 10'b0000100001;
    pxcRom[3659] <= 10'b0000010001;
    pxcRom[3660] <= 10'b0000001001;
    pxcRom[3661] <= 10'b0000000100;
    pxcRom[3662] <= 10'b0000000010;
    pxcRom[3663] <= 10'b0000000001;
    pxcRom[3664] <= 10'b0000000000;
    pxcRom[3665] <= 10'b0000000000;
    pxcRom[3666] <= 10'b0000000000;
    pxcRom[3667] <= 10'b0000000000;
    pxcRom[3668] <= 10'b0000000000;
    pxcRom[3669] <= 10'b0000000000;
    pxcRom[3670] <= 10'b0000000000;
    pxcRom[3671] <= 10'b0000000000;
    pxcRom[3672] <= 10'b0000000000;
    pxcRom[3673] <= 10'b0000000001;
    pxcRom[3674] <= 10'b0000000011;
    pxcRom[3675] <= 10'b0000000100;
    pxcRom[3676] <= 10'b0000000101;
    pxcRom[3677] <= 10'b0000000110;
    pxcRom[3678] <= 10'b0000000111;
    pxcRom[3679] <= 10'b0000001100;
    pxcRom[3680] <= 10'b0000010100;
    pxcRom[3681] <= 10'b0000100010;
    pxcRom[3682] <= 10'b0000110010;
    pxcRom[3683] <= 10'b0000111100;
    pxcRom[3684] <= 10'b0000111001;
    pxcRom[3685] <= 10'b0000101001;
    pxcRom[3686] <= 10'b0000011001;
    pxcRom[3687] <= 10'b0000001101;
    pxcRom[3688] <= 10'b0000000111;
    pxcRom[3689] <= 10'b0000000011;
    pxcRom[3690] <= 10'b0000000001;
    pxcRom[3691] <= 10'b0000000000;
    pxcRom[3692] <= 10'b0000000000;
    pxcRom[3693] <= 10'b0000000000;
    pxcRom[3694] <= 10'b0000000000;
    pxcRom[3695] <= 10'b0000000000;
    pxcRom[3696] <= 10'b0000000000;
    pxcRom[3697] <= 10'b0000000000;
    pxcRom[3698] <= 10'b0000000000;
    pxcRom[3699] <= 10'b0000000000;
    pxcRom[3700] <= 10'b0000000000;
    pxcRom[3701] <= 10'b0000000000;
    pxcRom[3702] <= 10'b0000000001;
    pxcRom[3703] <= 10'b0000000001;
    pxcRom[3704] <= 10'b0000000001;
    pxcRom[3705] <= 10'b0000000011;
    pxcRom[3706] <= 10'b0000000101;
    pxcRom[3707] <= 10'b0000001100;
    pxcRom[3708] <= 10'b0000010101;
    pxcRom[3709] <= 10'b0000100001;
    pxcRom[3710] <= 10'b0000101100;
    pxcRom[3711] <= 10'b0000110001;
    pxcRom[3712] <= 10'b0000101101;
    pxcRom[3713] <= 10'b0000100010;
    pxcRom[3714] <= 10'b0000010101;
    pxcRom[3715] <= 10'b0000001100;
    pxcRom[3716] <= 10'b0000000110;
    pxcRom[3717] <= 10'b0000000011;
    pxcRom[3718] <= 10'b0000000001;
    pxcRom[3719] <= 10'b0000000000;
    pxcRom[3720] <= 10'b0000000000;
    pxcRom[3721] <= 10'b0000000000;
    pxcRom[3722] <= 10'b0000000000;
    pxcRom[3723] <= 10'b0000000000;
    pxcRom[3724] <= 10'b0000000000;
    pxcRom[3725] <= 10'b0000000000;
    pxcRom[3726] <= 10'b0000000000;
    pxcRom[3727] <= 10'b0000000000;
    pxcRom[3728] <= 10'b0000000000;
    pxcRom[3729] <= 10'b0000000000;
    pxcRom[3730] <= 10'b0000000000;
    pxcRom[3731] <= 10'b0000000000;
    pxcRom[3732] <= 10'b0000000001;
    pxcRom[3733] <= 10'b0000000011;
    pxcRom[3734] <= 10'b0000001000;
    pxcRom[3735] <= 10'b0000001110;
    pxcRom[3736] <= 10'b0000010111;
    pxcRom[3737] <= 10'b0000100000;
    pxcRom[3738] <= 10'b0000100110;
    pxcRom[3739] <= 10'b0000101001;
    pxcRom[3740] <= 10'b0000100110;
    pxcRom[3741] <= 10'b0000011101;
    pxcRom[3742] <= 10'b0000010100;
    pxcRom[3743] <= 10'b0000001100;
    pxcRom[3744] <= 10'b0000000110;
    pxcRom[3745] <= 10'b0000000011;
    pxcRom[3746] <= 10'b0000000001;
    pxcRom[3747] <= 10'b0000000000;
    pxcRom[3748] <= 10'b0000000000;
    pxcRom[3749] <= 10'b0000000000;
    pxcRom[3750] <= 10'b0000000000;
    pxcRom[3751] <= 10'b0000000000;
    pxcRom[3752] <= 10'b0000000000;
    pxcRom[3753] <= 10'b0000000000;
    pxcRom[3754] <= 10'b0000000000;
    pxcRom[3755] <= 10'b0000000000;
    pxcRom[3756] <= 10'b0000000000;
    pxcRom[3757] <= 10'b0000000000;
    pxcRom[3758] <= 10'b0000000000;
    pxcRom[3759] <= 10'b0000000000;
    pxcRom[3760] <= 10'b0000000010;
    pxcRom[3761] <= 10'b0000000101;
    pxcRom[3762] <= 10'b0000001010;
    pxcRom[3763] <= 10'b0000010000;
    pxcRom[3764] <= 10'b0000011000;
    pxcRom[3765] <= 10'b0000011110;
    pxcRom[3766] <= 10'b0000100010;
    pxcRom[3767] <= 10'b0000100011;
    pxcRom[3768] <= 10'b0000100001;
    pxcRom[3769] <= 10'b0000011010;
    pxcRom[3770] <= 10'b0000010010;
    pxcRom[3771] <= 10'b0000001100;
    pxcRom[3772] <= 10'b0000000111;
    pxcRom[3773] <= 10'b0000000011;
    pxcRom[3774] <= 10'b0000000001;
    pxcRom[3775] <= 10'b0000000000;
    pxcRom[3776] <= 10'b0000000000;
    pxcRom[3777] <= 10'b0000000000;
    pxcRom[3778] <= 10'b0000000000;
    pxcRom[3779] <= 10'b0000000000;
    pxcRom[3780] <= 10'b0000000000;
    pxcRom[3781] <= 10'b0000000000;
    pxcRom[3782] <= 10'b0000000000;
    pxcRom[3783] <= 10'b0000000000;
    pxcRom[3784] <= 10'b0000000000;
    pxcRom[3785] <= 10'b0000000000;
    pxcRom[3786] <= 10'b0000000000;
    pxcRom[3787] <= 10'b0000000001;
    pxcRom[3788] <= 10'b0000000010;
    pxcRom[3789] <= 10'b0000000101;
    pxcRom[3790] <= 10'b0000001010;
    pxcRom[3791] <= 10'b0000010000;
    pxcRom[3792] <= 10'b0000010101;
    pxcRom[3793] <= 10'b0000011010;
    pxcRom[3794] <= 10'b0000011100;
    pxcRom[3795] <= 10'b0000011101;
    pxcRom[3796] <= 10'b0000011011;
    pxcRom[3797] <= 10'b0000010111;
    pxcRom[3798] <= 10'b0000010000;
    pxcRom[3799] <= 10'b0000001011;
    pxcRom[3800] <= 10'b0000000110;
    pxcRom[3801] <= 10'b0000000011;
    pxcRom[3802] <= 10'b0000000001;
    pxcRom[3803] <= 10'b0000000000;
    pxcRom[3804] <= 10'b0000000000;
    pxcRom[3805] <= 10'b0000000000;
    pxcRom[3806] <= 10'b0000000000;
    pxcRom[3807] <= 10'b0000000000;
    pxcRom[3808] <= 10'b0000000000;
    pxcRom[3809] <= 10'b0000000000;
    pxcRom[3810] <= 10'b0000000000;
    pxcRom[3811] <= 10'b0000000000;
    pxcRom[3812] <= 10'b0000000000;
    pxcRom[3813] <= 10'b0000000000;
    pxcRom[3814] <= 10'b0000000000;
    pxcRom[3815] <= 10'b0000000001;
    pxcRom[3816] <= 10'b0000000010;
    pxcRom[3817] <= 10'b0000000100;
    pxcRom[3818] <= 10'b0000000111;
    pxcRom[3819] <= 10'b0000001011;
    pxcRom[3820] <= 10'b0000001110;
    pxcRom[3821] <= 10'b0000010000;
    pxcRom[3822] <= 10'b0000010001;
    pxcRom[3823] <= 10'b0000010010;
    pxcRom[3824] <= 10'b0000010001;
    pxcRom[3825] <= 10'b0000001110;
    pxcRom[3826] <= 10'b0000001010;
    pxcRom[3827] <= 10'b0000000111;
    pxcRom[3828] <= 10'b0000000100;
    pxcRom[3829] <= 10'b0000000010;
    pxcRom[3830] <= 10'b0000000001;
    pxcRom[3831] <= 10'b0000000000;
    pxcRom[3832] <= 10'b0000000000;
    pxcRom[3833] <= 10'b0000000000;
    pxcRom[3834] <= 10'b0000000000;
    pxcRom[3835] <= 10'b0000000000;
    pxcRom[3836] <= 10'b0000000000;
    pxcRom[3837] <= 10'b0000000000;
    pxcRom[3838] <= 10'b0000000000;
    pxcRom[3839] <= 10'b0000000000;
    pxcRom[3840] <= 10'b0000000000;
    pxcRom[3841] <= 10'b0000000000;
    pxcRom[3842] <= 10'b0000000000;
    pxcRom[3843] <= 10'b0000000000;
    pxcRom[3844] <= 10'b0000000000;
    pxcRom[3845] <= 10'b0000000001;
    pxcRom[3846] <= 10'b0000000010;
    pxcRom[3847] <= 10'b0000000010;
    pxcRom[3848] <= 10'b0000000011;
    pxcRom[3849] <= 10'b0000000100;
    pxcRom[3850] <= 10'b0000000100;
    pxcRom[3851] <= 10'b0000000100;
    pxcRom[3852] <= 10'b0000000100;
    pxcRom[3853] <= 10'b0000000011;
    pxcRom[3854] <= 10'b0000000010;
    pxcRom[3855] <= 10'b0000000001;
    pxcRom[3856] <= 10'b0000000000;
    pxcRom[3857] <= 10'b0000000000;
    pxcRom[3858] <= 10'b0000000000;
    pxcRom[3859] <= 10'b0000000000;
    pxcRom[3860] <= 10'b0000000000;
    pxcRom[3861] <= 10'b0000000000;
    pxcRom[3862] <= 10'b0000000000;
    pxcRom[3863] <= 10'b0000000000;
    pxcRom[3864] <= 10'b0000000000;
    pxcRom[3865] <= 10'b0000000000;
    pxcRom[3866] <= 10'b0000000000;
    pxcRom[3867] <= 10'b0000000000;
    pxcRom[3868] <= 10'b0000000000;
    pxcRom[3869] <= 10'b0000000000;
    pxcRom[3870] <= 10'b0000000000;
    pxcRom[3871] <= 10'b0000000000;
    pxcRom[3872] <= 10'b0000000000;
    pxcRom[3873] <= 10'b0000000000;
    pxcRom[3874] <= 10'b0000000000;
    pxcRom[3875] <= 10'b0000000000;
    pxcRom[3876] <= 10'b0000000000;
    pxcRom[3877] <= 10'b0000000000;
    pxcRom[3878] <= 10'b0000000000;
    pxcRom[3879] <= 10'b0000000000;
    pxcRom[3880] <= 10'b0000000000;
    pxcRom[3881] <= 10'b0000000000;
    pxcRom[3882] <= 10'b0000000000;
    pxcRom[3883] <= 10'b0000000000;
    pxcRom[3884] <= 10'b0000000000;
    pxcRom[3885] <= 10'b0000000000;
    pxcRom[3886] <= 10'b0000000000;
    pxcRom[3887] <= 10'b0000000000;
    pxcRom[3888] <= 10'b0000000000;
    pxcRom[3889] <= 10'b0000000000;
    pxcRom[3890] <= 10'b0000000000;
    pxcRom[3891] <= 10'b0000000000;
    pxcRom[3892] <= 10'b0000000000;
    pxcRom[3893] <= 10'b0000000000;
    pxcRom[3894] <= 10'b0000000000;
    pxcRom[3895] <= 10'b0000000000;
    pxcRom[3896] <= 10'b0000000000;
    pxcRom[3897] <= 10'b0000000000;
    pxcRom[3898] <= 10'b0000000000;
    pxcRom[3899] <= 10'b0000000000;
    pxcRom[3900] <= 10'b0000000000;
    pxcRom[3901] <= 10'b0000000000;
    pxcRom[3902] <= 10'b0000000000;
    pxcRom[3903] <= 10'b0000000000;
    pxcRom[3904] <= 10'b0000000000;
    pxcRom[3905] <= 10'b0000000000;
    pxcRom[3906] <= 10'b0000000000;
    pxcRom[3907] <= 10'b0000000000;
    pxcRom[3908] <= 10'b0000000000;
    pxcRom[3909] <= 10'b0000000000;
    pxcRom[3910] <= 10'b0000000000;
    pxcRom[3911] <= 10'b0000000000;
    pxcRom[3912] <= 10'b0000000000;
    pxcRom[3913] <= 10'b0000000000;
    pxcRom[3914] <= 10'b0000000000;
    pxcRom[3915] <= 10'b0000000000;
    pxcRom[3916] <= 10'b0000000000;
    pxcRom[3917] <= 10'b0000000000;
    pxcRom[3918] <= 10'b0000000000;
    pxcRom[3919] <= 10'b0000000000;
    pxcRom[3920] <= 10'b0000000000;
    pxcRom[3921] <= 10'b0000000000;
    pxcRom[3922] <= 10'b0000000000;
    pxcRom[3923] <= 10'b0000000000;
    pxcRom[3924] <= 10'b0000000000;
    pxcRom[3925] <= 10'b0000000000;
    pxcRom[3926] <= 10'b0000000000;
    pxcRom[3927] <= 10'b0000000000;
    pxcRom[3928] <= 10'b0000000000;
    pxcRom[3929] <= 10'b0000000000;
    pxcRom[3930] <= 10'b0000000000;
    pxcRom[3931] <= 10'b0000000000;
    pxcRom[3932] <= 10'b0000000000;
    pxcRom[3933] <= 10'b0000000000;
    pxcRom[3934] <= 10'b0000000000;
    pxcRom[3935] <= 10'b0000000000;
    pxcRom[3936] <= 10'b0000000000;
    pxcRom[3937] <= 10'b0000000000;
    pxcRom[3938] <= 10'b0000000000;
    pxcRom[3939] <= 10'b0000000000;
    pxcRom[3940] <= 10'b0000000000;
    pxcRom[3941] <= 10'b0000000000;
    pxcRom[3942] <= 10'b0000000000;
    pxcRom[3943] <= 10'b0000000000;
    pxcRom[3944] <= 10'b0000000000;
    pxcRom[3945] <= 10'b0000000000;
    pxcRom[3946] <= 10'b0000000000;
    pxcRom[3947] <= 10'b0000000000;
    pxcRom[3948] <= 10'b0000000000;
    pxcRom[3949] <= 10'b0000000000;
    pxcRom[3950] <= 10'b0000000000;
    pxcRom[3951] <= 10'b0000000000;
    pxcRom[3952] <= 10'b0000000000;
    pxcRom[3953] <= 10'b0000000000;
    pxcRom[3954] <= 10'b0000000000;
    pxcRom[3955] <= 10'b0000000000;
    pxcRom[3956] <= 10'b0000000000;
    pxcRom[3957] <= 10'b0000000000;
    pxcRom[3958] <= 10'b0000000000;
    pxcRom[3959] <= 10'b0000000000;
    pxcRom[3960] <= 10'b0000000000;
    pxcRom[3961] <= 10'b0000000000;
    pxcRom[3962] <= 10'b0000000000;
    pxcRom[3963] <= 10'b0000000000;
    pxcRom[3964] <= 10'b0000000000;
    pxcRom[3965] <= 10'b0000000000;
    pxcRom[3966] <= 10'b0000000000;
    pxcRom[3967] <= 10'b0000000000;
    pxcRom[3968] <= 10'b0000000000;
    pxcRom[3969] <= 10'b0000000000;
    pxcRom[3970] <= 10'b0000000000;
    pxcRom[3971] <= 10'b0000000000;
    pxcRom[3972] <= 10'b0000000000;
    pxcRom[3973] <= 10'b0000000000;
    pxcRom[3974] <= 10'b0000000000;
    pxcRom[3975] <= 10'b0000000000;
    pxcRom[3976] <= 10'b0000000000;
    pxcRom[3977] <= 10'b0000000000;
    pxcRom[3978] <= 10'b0000000000;
    pxcRom[3979] <= 10'b0000000000;
    pxcRom[3980] <= 10'b0000000000;
    pxcRom[3981] <= 10'b0000000000;
    pxcRom[3982] <= 10'b0000000000;
    pxcRom[3983] <= 10'b0000000000;
    pxcRom[3984] <= 10'b0000000000;
    pxcRom[3985] <= 10'b0000000000;
    pxcRom[3986] <= 10'b0000000000;
    pxcRom[3987] <= 10'b0000000000;
    pxcRom[3988] <= 10'b0000000000;
    pxcRom[3989] <= 10'b0000000000;
    pxcRom[3990] <= 10'b0000000000;
    pxcRom[3991] <= 10'b0000000000;
    pxcRom[3992] <= 10'b0000000000;
    pxcRom[3993] <= 10'b0000000000;
    pxcRom[3994] <= 10'b0000000000;
    pxcRom[3995] <= 10'b0000000000;
    pxcRom[3996] <= 10'b0000000000;
    pxcRom[3997] <= 10'b0000000000;
    pxcRom[3998] <= 10'b0000000000;
    pxcRom[3999] <= 10'b0000000000;
    pxcRom[4000] <= 10'b0000000000;
    pxcRom[4001] <= 10'b0000000000;
    pxcRom[4002] <= 10'b0000000000;
    pxcRom[4003] <= 10'b0000000000;
    pxcRom[4004] <= 10'b0000000000;
    pxcRom[4005] <= 10'b0000000000;
    pxcRom[4006] <= 10'b0000000000;
    pxcRom[4007] <= 10'b0000000000;
    pxcRom[4008] <= 10'b0000000000;
    pxcRom[4009] <= 10'b0000000000;
    pxcRom[4010] <= 10'b0000000000;
    pxcRom[4011] <= 10'b0000000000;
    pxcRom[4012] <= 10'b0000000000;
    pxcRom[4013] <= 10'b0000000000;
    pxcRom[4014] <= 10'b0000000000;
    pxcRom[4015] <= 10'b0000000000;
    pxcRom[4016] <= 10'b0000000000;
    pxcRom[4017] <= 10'b0000000000;
    pxcRom[4018] <= 10'b0000000000;
    pxcRom[4019] <= 10'b0000000001;
    pxcRom[4020] <= 10'b0000000001;
    pxcRom[4021] <= 10'b0000000001;
    pxcRom[4022] <= 10'b0000000001;
    pxcRom[4023] <= 10'b0000000001;
    pxcRom[4024] <= 10'b0000000000;
    pxcRom[4025] <= 10'b0000000000;
    pxcRom[4026] <= 10'b0000000000;
    pxcRom[4027] <= 10'b0000000000;
    pxcRom[4028] <= 10'b0000000000;
    pxcRom[4029] <= 10'b0000000000;
    pxcRom[4030] <= 10'b0000000000;
    pxcRom[4031] <= 10'b0000000000;
    pxcRom[4032] <= 10'b0000000000;
    pxcRom[4033] <= 10'b0000000000;
    pxcRom[4034] <= 10'b0000000000;
    pxcRom[4035] <= 10'b0000000000;
    pxcRom[4036] <= 10'b0000000000;
    pxcRom[4037] <= 10'b0000000000;
    pxcRom[4038] <= 10'b0000000000;
    pxcRom[4039] <= 10'b0000000000;
    pxcRom[4040] <= 10'b0000000000;
    pxcRom[4041] <= 10'b0000000001;
    pxcRom[4042] <= 10'b0000000010;
    pxcRom[4043] <= 10'b0000000100;
    pxcRom[4044] <= 10'b0000000101;
    pxcRom[4045] <= 10'b0000000111;
    pxcRom[4046] <= 10'b0000001000;
    pxcRom[4047] <= 10'b0000001001;
    pxcRom[4048] <= 10'b0000001011;
    pxcRom[4049] <= 10'b0000001011;
    pxcRom[4050] <= 10'b0000001010;
    pxcRom[4051] <= 10'b0000001001;
    pxcRom[4052] <= 10'b0000001000;
    pxcRom[4053] <= 10'b0000000111;
    pxcRom[4054] <= 10'b0000000101;
    pxcRom[4055] <= 10'b0000000100;
    pxcRom[4056] <= 10'b0000000010;
    pxcRom[4057] <= 10'b0000000000;
    pxcRom[4058] <= 10'b0000000000;
    pxcRom[4059] <= 10'b0000000000;
    pxcRom[4060] <= 10'b0000000000;
    pxcRom[4061] <= 10'b0000000000;
    pxcRom[4062] <= 10'b0000000000;
    pxcRom[4063] <= 10'b0000000000;
    pxcRom[4064] <= 10'b0000000000;
    pxcRom[4065] <= 10'b0000000000;
    pxcRom[4066] <= 10'b0000000000;
    pxcRom[4067] <= 10'b0000000001;
    pxcRom[4068] <= 10'b0000000011;
    pxcRom[4069] <= 10'b0000000110;
    pxcRom[4070] <= 10'b0000001010;
    pxcRom[4071] <= 10'b0000001111;
    pxcRom[4072] <= 10'b0000010101;
    pxcRom[4073] <= 10'b0000011010;
    pxcRom[4074] <= 10'b0000011111;
    pxcRom[4075] <= 10'b0000100010;
    pxcRom[4076] <= 10'b0000100100;
    pxcRom[4077] <= 10'b0000100100;
    pxcRom[4078] <= 10'b0000100011;
    pxcRom[4079] <= 10'b0000100000;
    pxcRom[4080] <= 10'b0000011100;
    pxcRom[4081] <= 10'b0000010111;
    pxcRom[4082] <= 10'b0000010011;
    pxcRom[4083] <= 10'b0000001101;
    pxcRom[4084] <= 10'b0000001000;
    pxcRom[4085] <= 10'b0000000011;
    pxcRom[4086] <= 10'b0000000000;
    pxcRom[4087] <= 10'b0000000000;
    pxcRom[4088] <= 10'b0000000000;
    pxcRom[4089] <= 10'b0000000000;
    pxcRom[4090] <= 10'b0000000000;
    pxcRom[4091] <= 10'b0000000000;
    pxcRom[4092] <= 10'b0000000000;
    pxcRom[4093] <= 10'b0000000000;
    pxcRom[4094] <= 10'b0000000001;
    pxcRom[4095] <= 10'b0000000011;
    pxcRom[4096] <= 10'b0000000110;
    pxcRom[4097] <= 10'b0000001100;
    pxcRom[4098] <= 10'b0000010100;
    pxcRom[4099] <= 10'b0000011110;
    pxcRom[4100] <= 10'b0000101001;
    pxcRom[4101] <= 10'b0000110010;
    pxcRom[4102] <= 10'b0000111001;
    pxcRom[4103] <= 10'b0000111101;
    pxcRom[4104] <= 10'b0000111101;
    pxcRom[4105] <= 10'b0000111110;
    pxcRom[4106] <= 10'b0000111010;
    pxcRom[4107] <= 10'b0000110101;
    pxcRom[4108] <= 10'b0000101110;
    pxcRom[4109] <= 10'b0000100110;
    pxcRom[4110] <= 10'b0000011111;
    pxcRom[4111] <= 10'b0000011000;
    pxcRom[4112] <= 10'b0000001111;
    pxcRom[4113] <= 10'b0000000110;
    pxcRom[4114] <= 10'b0000000001;
    pxcRom[4115] <= 10'b0000000000;
    pxcRom[4116] <= 10'b0000000000;
    pxcRom[4117] <= 10'b0000000000;
    pxcRom[4118] <= 10'b0000000000;
    pxcRom[4119] <= 10'b0000000000;
    pxcRom[4120] <= 10'b0000000000;
    pxcRom[4121] <= 10'b0000000000;
    pxcRom[4122] <= 10'b0000000010;
    pxcRom[4123] <= 10'b0000000101;
    pxcRom[4124] <= 10'b0000001010;
    pxcRom[4125] <= 10'b0000010011;
    pxcRom[4126] <= 10'b0000011111;
    pxcRom[4127] <= 10'b0000101101;
    pxcRom[4128] <= 10'b0000111011;
    pxcRom[4129] <= 10'b0001000100;
    pxcRom[4130] <= 10'b0001001000;
    pxcRom[4131] <= 10'b0001001001;
    pxcRom[4132] <= 10'b0001000111;
    pxcRom[4133] <= 10'b0001000100;
    pxcRom[4134] <= 10'b0001000000;
    pxcRom[4135] <= 10'b0000111010;
    pxcRom[4136] <= 10'b0000110011;
    pxcRom[4137] <= 10'b0000101011;
    pxcRom[4138] <= 10'b0000100011;
    pxcRom[4139] <= 10'b0000011100;
    pxcRom[4140] <= 10'b0000010011;
    pxcRom[4141] <= 10'b0000001001;
    pxcRom[4142] <= 10'b0000000001;
    pxcRom[4143] <= 10'b0000000000;
    pxcRom[4144] <= 10'b0000000000;
    pxcRom[4145] <= 10'b0000000000;
    pxcRom[4146] <= 10'b0000000000;
    pxcRom[4147] <= 10'b0000000000;
    pxcRom[4148] <= 10'b0000000000;
    pxcRom[4149] <= 10'b0000000001;
    pxcRom[4150] <= 10'b0000000011;
    pxcRom[4151] <= 10'b0000000111;
    pxcRom[4152] <= 10'b0000001111;
    pxcRom[4153] <= 10'b0000011010;
    pxcRom[4154] <= 10'b0000101001;
    pxcRom[4155] <= 10'b0000111010;
    pxcRom[4156] <= 10'b0001000011;
    pxcRom[4157] <= 10'b0001000110;
    pxcRom[4158] <= 10'b0001000011;
    pxcRom[4159] <= 10'b0000111111;
    pxcRom[4160] <= 10'b0000111010;
    pxcRom[4161] <= 10'b0000110110;
    pxcRom[4162] <= 10'b0000110000;
    pxcRom[4163] <= 10'b0000101011;
    pxcRom[4164] <= 10'b0000100110;
    pxcRom[4165] <= 10'b0000100010;
    pxcRom[4166] <= 10'b0000011100;
    pxcRom[4167] <= 10'b0000010111;
    pxcRom[4168] <= 10'b0000010001;
    pxcRom[4169] <= 10'b0000001000;
    pxcRom[4170] <= 10'b0000000001;
    pxcRom[4171] <= 10'b0000000000;
    pxcRom[4172] <= 10'b0000000000;
    pxcRom[4173] <= 10'b0000000000;
    pxcRom[4174] <= 10'b0000000000;
    pxcRom[4175] <= 10'b0000000000;
    pxcRom[4176] <= 10'b0000000000;
    pxcRom[4177] <= 10'b0000000001;
    pxcRom[4178] <= 10'b0000000100;
    pxcRom[4179] <= 10'b0000001001;
    pxcRom[4180] <= 10'b0000010011;
    pxcRom[4181] <= 10'b0000100001;
    pxcRom[4182] <= 10'b0000110011;
    pxcRom[4183] <= 10'b0001000011;
    pxcRom[4184] <= 10'b0001000101;
    pxcRom[4185] <= 10'b0000111101;
    pxcRom[4186] <= 10'b0000110011;
    pxcRom[4187] <= 10'b0000101011;
    pxcRom[4188] <= 10'b0000100101;
    pxcRom[4189] <= 10'b0000100001;
    pxcRom[4190] <= 10'b0000011101;
    pxcRom[4191] <= 10'b0000011010;
    pxcRom[4192] <= 10'b0000010111;
    pxcRom[4193] <= 10'b0000010100;
    pxcRom[4194] <= 10'b0000010001;
    pxcRom[4195] <= 10'b0000001111;
    pxcRom[4196] <= 10'b0000001011;
    pxcRom[4197] <= 10'b0000000101;
    pxcRom[4198] <= 10'b0000000001;
    pxcRom[4199] <= 10'b0000000000;
    pxcRom[4200] <= 10'b0000000000;
    pxcRom[4201] <= 10'b0000000000;
    pxcRom[4202] <= 10'b0000000000;
    pxcRom[4203] <= 10'b0000000000;
    pxcRom[4204] <= 10'b0000000000;
    pxcRom[4205] <= 10'b0000000001;
    pxcRom[4206] <= 10'b0000000101;
    pxcRom[4207] <= 10'b0000001100;
    pxcRom[4208] <= 10'b0000011000;
    pxcRom[4209] <= 10'b0000101100;
    pxcRom[4210] <= 10'b0001000001;
    pxcRom[4211] <= 10'b0001001101;
    pxcRom[4212] <= 10'b0001001000;
    pxcRom[4213] <= 10'b0000111000;
    pxcRom[4214] <= 10'b0000101001;
    pxcRom[4215] <= 10'b0000100000;
    pxcRom[4216] <= 10'b0000011001;
    pxcRom[4217] <= 10'b0000010011;
    pxcRom[4218] <= 10'b0000010000;
    pxcRom[4219] <= 10'b0000001101;
    pxcRom[4220] <= 10'b0000001011;
    pxcRom[4221] <= 10'b0000001001;
    pxcRom[4222] <= 10'b0000000111;
    pxcRom[4223] <= 10'b0000000110;
    pxcRom[4224] <= 10'b0000000101;
    pxcRom[4225] <= 10'b0000000010;
    pxcRom[4226] <= 10'b0000000000;
    pxcRom[4227] <= 10'b0000000000;
    pxcRom[4228] <= 10'b0000000000;
    pxcRom[4229] <= 10'b0000000000;
    pxcRom[4230] <= 10'b0000000000;
    pxcRom[4231] <= 10'b0000000000;
    pxcRom[4232] <= 10'b0000000000;
    pxcRom[4233] <= 10'b0000000010;
    pxcRom[4234] <= 10'b0000000110;
    pxcRom[4235] <= 10'b0000001111;
    pxcRom[4236] <= 10'b0000011111;
    pxcRom[4237] <= 10'b0000110110;
    pxcRom[4238] <= 10'b0001010010;
    pxcRom[4239] <= 10'b0001011101;
    pxcRom[4240] <= 10'b0001001110;
    pxcRom[4241] <= 10'b0000111000;
    pxcRom[4242] <= 10'b0000101000;
    pxcRom[4243] <= 10'b0000011110;
    pxcRom[4244] <= 10'b0000010111;
    pxcRom[4245] <= 10'b0000010001;
    pxcRom[4246] <= 10'b0000001100;
    pxcRom[4247] <= 10'b0000001000;
    pxcRom[4248] <= 10'b0000000101;
    pxcRom[4249] <= 10'b0000000011;
    pxcRom[4250] <= 10'b0000000010;
    pxcRom[4251] <= 10'b0000000010;
    pxcRom[4252] <= 10'b0000000001;
    pxcRom[4253] <= 10'b0000000000;
    pxcRom[4254] <= 10'b0000000000;
    pxcRom[4255] <= 10'b0000000000;
    pxcRom[4256] <= 10'b0000000000;
    pxcRom[4257] <= 10'b0000000000;
    pxcRom[4258] <= 10'b0000000000;
    pxcRom[4259] <= 10'b0000000000;
    pxcRom[4260] <= 10'b0000000000;
    pxcRom[4261] <= 10'b0000000010;
    pxcRom[4262] <= 10'b0000000111;
    pxcRom[4263] <= 10'b0000010001;
    pxcRom[4264] <= 10'b0000100100;
    pxcRom[4265] <= 10'b0001000011;
    pxcRom[4266] <= 10'b0001100101;
    pxcRom[4267] <= 10'b0001101110;
    pxcRom[4268] <= 10'b0001011000;
    pxcRom[4269] <= 10'b0001000001;
    pxcRom[4270] <= 10'b0000110001;
    pxcRom[4271] <= 10'b0000100111;
    pxcRom[4272] <= 10'b0000011111;
    pxcRom[4273] <= 10'b0000011000;
    pxcRom[4274] <= 10'b0000010000;
    pxcRom[4275] <= 10'b0000001001;
    pxcRom[4276] <= 10'b0000000101;
    pxcRom[4277] <= 10'b0000000010;
    pxcRom[4278] <= 10'b0000000001;
    pxcRom[4279] <= 10'b0000000000;
    pxcRom[4280] <= 10'b0000000000;
    pxcRom[4281] <= 10'b0000000000;
    pxcRom[4282] <= 10'b0000000000;
    pxcRom[4283] <= 10'b0000000000;
    pxcRom[4284] <= 10'b0000000000;
    pxcRom[4285] <= 10'b0000000000;
    pxcRom[4286] <= 10'b0000000000;
    pxcRom[4287] <= 10'b0000000000;
    pxcRom[4288] <= 10'b0000000000;
    pxcRom[4289] <= 10'b0000000010;
    pxcRom[4290] <= 10'b0000000111;
    pxcRom[4291] <= 10'b0000010010;
    pxcRom[4292] <= 10'b0000100110;
    pxcRom[4293] <= 10'b0001000110;
    pxcRom[4294] <= 10'b0001100110;
    pxcRom[4295] <= 10'b0001101100;
    pxcRom[4296] <= 10'b0001011101;
    pxcRom[4297] <= 10'b0001001100;
    pxcRom[4298] <= 10'b0000111111;
    pxcRom[4299] <= 10'b0000110101;
    pxcRom[4300] <= 10'b0000101011;
    pxcRom[4301] <= 10'b0000100010;
    pxcRom[4302] <= 10'b0000011010;
    pxcRom[4303] <= 10'b0000010000;
    pxcRom[4304] <= 10'b0000001001;
    pxcRom[4305] <= 10'b0000000100;
    pxcRom[4306] <= 10'b0000000001;
    pxcRom[4307] <= 10'b0000000000;
    pxcRom[4308] <= 10'b0000000000;
    pxcRom[4309] <= 10'b0000000000;
    pxcRom[4310] <= 10'b0000000000;
    pxcRom[4311] <= 10'b0000000000;
    pxcRom[4312] <= 10'b0000000000;
    pxcRom[4313] <= 10'b0000000000;
    pxcRom[4314] <= 10'b0000000000;
    pxcRom[4315] <= 10'b0000000000;
    pxcRom[4316] <= 10'b0000000000;
    pxcRom[4317] <= 10'b0000000010;
    pxcRom[4318] <= 10'b0000000110;
    pxcRom[4319] <= 10'b0000001111;
    pxcRom[4320] <= 10'b0000100000;
    pxcRom[4321] <= 10'b0000111000;
    pxcRom[4322] <= 10'b0001001011;
    pxcRom[4323] <= 10'b0001010001;
    pxcRom[4324] <= 10'b0001001100;
    pxcRom[4325] <= 10'b0001000011;
    pxcRom[4326] <= 10'b0000111101;
    pxcRom[4327] <= 10'b0000110111;
    pxcRom[4328] <= 10'b0000110010;
    pxcRom[4329] <= 10'b0000101100;
    pxcRom[4330] <= 10'b0000100011;
    pxcRom[4331] <= 10'b0000011000;
    pxcRom[4332] <= 10'b0000001110;
    pxcRom[4333] <= 10'b0000000111;
    pxcRom[4334] <= 10'b0000000011;
    pxcRom[4335] <= 10'b0000000001;
    pxcRom[4336] <= 10'b0000000000;
    pxcRom[4337] <= 10'b0000000000;
    pxcRom[4338] <= 10'b0000000000;
    pxcRom[4339] <= 10'b0000000000;
    pxcRom[4340] <= 10'b0000000000;
    pxcRom[4341] <= 10'b0000000000;
    pxcRom[4342] <= 10'b0000000000;
    pxcRom[4343] <= 10'b0000000000;
    pxcRom[4344] <= 10'b0000000000;
    pxcRom[4345] <= 10'b0000000010;
    pxcRom[4346] <= 10'b0000000101;
    pxcRom[4347] <= 10'b0000001011;
    pxcRom[4348] <= 10'b0000010110;
    pxcRom[4349] <= 10'b0000100010;
    pxcRom[4350] <= 10'b0000101011;
    pxcRom[4351] <= 10'b0000101110;
    pxcRom[4352] <= 10'b0000101101;
    pxcRom[4353] <= 10'b0000101101;
    pxcRom[4354] <= 10'b0000101101;
    pxcRom[4355] <= 10'b0000101110;
    pxcRom[4356] <= 10'b0000110000;
    pxcRom[4357] <= 10'b0000101110;
    pxcRom[4358] <= 10'b0000101010;
    pxcRom[4359] <= 10'b0000011111;
    pxcRom[4360] <= 10'b0000010011;
    pxcRom[4361] <= 10'b0000001010;
    pxcRom[4362] <= 10'b0000000101;
    pxcRom[4363] <= 10'b0000000010;
    pxcRom[4364] <= 10'b0000000000;
    pxcRom[4365] <= 10'b0000000000;
    pxcRom[4366] <= 10'b0000000000;
    pxcRom[4367] <= 10'b0000000000;
    pxcRom[4368] <= 10'b0000000000;
    pxcRom[4369] <= 10'b0000000000;
    pxcRom[4370] <= 10'b0000000000;
    pxcRom[4371] <= 10'b0000000000;
    pxcRom[4372] <= 10'b0000000000;
    pxcRom[4373] <= 10'b0000000010;
    pxcRom[4374] <= 10'b0000000101;
    pxcRom[4375] <= 10'b0000001000;
    pxcRom[4376] <= 10'b0000001101;
    pxcRom[4377] <= 10'b0000010010;
    pxcRom[4378] <= 10'b0000010101;
    pxcRom[4379] <= 10'b0000010110;
    pxcRom[4380] <= 10'b0000010111;
    pxcRom[4381] <= 10'b0000011001;
    pxcRom[4382] <= 10'b0000011101;
    pxcRom[4383] <= 10'b0000100011;
    pxcRom[4384] <= 10'b0000101010;
    pxcRom[4385] <= 10'b0000101111;
    pxcRom[4386] <= 10'b0000101101;
    pxcRom[4387] <= 10'b0000100011;
    pxcRom[4388] <= 10'b0000010111;
    pxcRom[4389] <= 10'b0000001101;
    pxcRom[4390] <= 10'b0000000110;
    pxcRom[4391] <= 10'b0000000010;
    pxcRom[4392] <= 10'b0000000000;
    pxcRom[4393] <= 10'b0000000000;
    pxcRom[4394] <= 10'b0000000000;
    pxcRom[4395] <= 10'b0000000000;
    pxcRom[4396] <= 10'b0000000000;
    pxcRom[4397] <= 10'b0000000000;
    pxcRom[4398] <= 10'b0000000000;
    pxcRom[4399] <= 10'b0000000000;
    pxcRom[4400] <= 10'b0000000001;
    pxcRom[4401] <= 10'b0000000101;
    pxcRom[4402] <= 10'b0000001001;
    pxcRom[4403] <= 10'b0000001011;
    pxcRom[4404] <= 10'b0000001010;
    pxcRom[4405] <= 10'b0000001010;
    pxcRom[4406] <= 10'b0000001010;
    pxcRom[4407] <= 10'b0000001011;
    pxcRom[4408] <= 10'b0000001011;
    pxcRom[4409] <= 10'b0000001111;
    pxcRom[4410] <= 10'b0000010110;
    pxcRom[4411] <= 10'b0000011110;
    pxcRom[4412] <= 10'b0000101000;
    pxcRom[4413] <= 10'b0000101111;
    pxcRom[4414] <= 10'b0000101110;
    pxcRom[4415] <= 10'b0000100101;
    pxcRom[4416] <= 10'b0000011000;
    pxcRom[4417] <= 10'b0000001110;
    pxcRom[4418] <= 10'b0000000111;
    pxcRom[4419] <= 10'b0000000011;
    pxcRom[4420] <= 10'b0000000001;
    pxcRom[4421] <= 10'b0000000000;
    pxcRom[4422] <= 10'b0000000000;
    pxcRom[4423] <= 10'b0000000000;
    pxcRom[4424] <= 10'b0000000000;
    pxcRom[4425] <= 10'b0000000000;
    pxcRom[4426] <= 10'b0000000000;
    pxcRom[4427] <= 10'b0000000000;
    pxcRom[4428] <= 10'b0000000010;
    pxcRom[4429] <= 10'b0000001000;
    pxcRom[4430] <= 10'b0000010000;
    pxcRom[4431] <= 10'b0000010001;
    pxcRom[4432] <= 10'b0000001111;
    pxcRom[4433] <= 10'b0000001100;
    pxcRom[4434] <= 10'b0000001010;
    pxcRom[4435] <= 10'b0000001001;
    pxcRom[4436] <= 10'b0000001010;
    pxcRom[4437] <= 10'b0000001110;
    pxcRom[4438] <= 10'b0000010110;
    pxcRom[4439] <= 10'b0000100000;
    pxcRom[4440] <= 10'b0000101010;
    pxcRom[4441] <= 10'b0000110001;
    pxcRom[4442] <= 10'b0000101111;
    pxcRom[4443] <= 10'b0000100100;
    pxcRom[4444] <= 10'b0000011000;
    pxcRom[4445] <= 10'b0000001110;
    pxcRom[4446] <= 10'b0000000111;
    pxcRom[4447] <= 10'b0000000011;
    pxcRom[4448] <= 10'b0000000001;
    pxcRom[4449] <= 10'b0000000000;
    pxcRom[4450] <= 10'b0000000000;
    pxcRom[4451] <= 10'b0000000000;
    pxcRom[4452] <= 10'b0000000000;
    pxcRom[4453] <= 10'b0000000000;
    pxcRom[4454] <= 10'b0000000000;
    pxcRom[4455] <= 10'b0000000000;
    pxcRom[4456] <= 10'b0000000011;
    pxcRom[4457] <= 10'b0000001011;
    pxcRom[4458] <= 10'b0000010111;
    pxcRom[4459] <= 10'b0000011101;
    pxcRom[4460] <= 10'b0000011100;
    pxcRom[4461] <= 10'b0000010111;
    pxcRom[4462] <= 10'b0000010011;
    pxcRom[4463] <= 10'b0000010000;
    pxcRom[4464] <= 10'b0000010001;
    pxcRom[4465] <= 10'b0000010101;
    pxcRom[4466] <= 10'b0000011101;
    pxcRom[4467] <= 10'b0000101000;
    pxcRom[4468] <= 10'b0000110001;
    pxcRom[4469] <= 10'b0000110100;
    pxcRom[4470] <= 10'b0000110000;
    pxcRom[4471] <= 10'b0000100011;
    pxcRom[4472] <= 10'b0000010111;
    pxcRom[4473] <= 10'b0000001101;
    pxcRom[4474] <= 10'b0000000111;
    pxcRom[4475] <= 10'b0000000011;
    pxcRom[4476] <= 10'b0000000000;
    pxcRom[4477] <= 10'b0000000000;
    pxcRom[4478] <= 10'b0000000000;
    pxcRom[4479] <= 10'b0000000000;
    pxcRom[4480] <= 10'b0000000000;
    pxcRom[4481] <= 10'b0000000000;
    pxcRom[4482] <= 10'b0000000000;
    pxcRom[4483] <= 10'b0000000000;
    pxcRom[4484] <= 10'b0000000010;
    pxcRom[4485] <= 10'b0000001011;
    pxcRom[4486] <= 10'b0000011010;
    pxcRom[4487] <= 10'b0000100110;
    pxcRom[4488] <= 10'b0000101100;
    pxcRom[4489] <= 10'b0000101100;
    pxcRom[4490] <= 10'b0000100111;
    pxcRom[4491] <= 10'b0000100011;
    pxcRom[4492] <= 10'b0000100010;
    pxcRom[4493] <= 10'b0000100110;
    pxcRom[4494] <= 10'b0000101101;
    pxcRom[4495] <= 10'b0000110110;
    pxcRom[4496] <= 10'b0000111011;
    pxcRom[4497] <= 10'b0000111001;
    pxcRom[4498] <= 10'b0000101110;
    pxcRom[4499] <= 10'b0000100000;
    pxcRom[4500] <= 10'b0000010100;
    pxcRom[4501] <= 10'b0000001011;
    pxcRom[4502] <= 10'b0000000101;
    pxcRom[4503] <= 10'b0000000010;
    pxcRom[4504] <= 10'b0000000000;
    pxcRom[4505] <= 10'b0000000000;
    pxcRom[4506] <= 10'b0000000000;
    pxcRom[4507] <= 10'b0000000000;
    pxcRom[4508] <= 10'b0000000000;
    pxcRom[4509] <= 10'b0000000000;
    pxcRom[4510] <= 10'b0000000000;
    pxcRom[4511] <= 10'b0000000000;
    pxcRom[4512] <= 10'b0000000010;
    pxcRom[4513] <= 10'b0000001000;
    pxcRom[4514] <= 10'b0000010110;
    pxcRom[4515] <= 10'b0000100111;
    pxcRom[4516] <= 10'b0000110110;
    pxcRom[4517] <= 10'b0000111111;
    pxcRom[4518] <= 10'b0001000010;
    pxcRom[4519] <= 10'b0001000000;
    pxcRom[4520] <= 10'b0001000000;
    pxcRom[4521] <= 10'b0001000001;
    pxcRom[4522] <= 10'b0001000110;
    pxcRom[4523] <= 10'b0001000111;
    pxcRom[4524] <= 10'b0001000100;
    pxcRom[4525] <= 10'b0000111000;
    pxcRom[4526] <= 10'b0000100111;
    pxcRom[4527] <= 10'b0000011001;
    pxcRom[4528] <= 10'b0000001110;
    pxcRom[4529] <= 10'b0000001000;
    pxcRom[4530] <= 10'b0000000011;
    pxcRom[4531] <= 10'b0000000001;
    pxcRom[4532] <= 10'b0000000000;
    pxcRom[4533] <= 10'b0000000000;
    pxcRom[4534] <= 10'b0000000000;
    pxcRom[4535] <= 10'b0000000000;
    pxcRom[4536] <= 10'b0000000000;
    pxcRom[4537] <= 10'b0000000000;
    pxcRom[4538] <= 10'b0000000000;
    pxcRom[4539] <= 10'b0000000000;
    pxcRom[4540] <= 10'b0000000001;
    pxcRom[4541] <= 10'b0000000100;
    pxcRom[4542] <= 10'b0000001110;
    pxcRom[4543] <= 10'b0000011100;
    pxcRom[4544] <= 10'b0000101110;
    pxcRom[4545] <= 10'b0001000000;
    pxcRom[4546] <= 10'b0001001101;
    pxcRom[4547] <= 10'b0001010101;
    pxcRom[4548] <= 10'b0001011000;
    pxcRom[4549] <= 10'b0001010110;
    pxcRom[4550] <= 10'b0001001111;
    pxcRom[4551] <= 10'b0001001000;
    pxcRom[4552] <= 10'b0000111011;
    pxcRom[4553] <= 10'b0000101011;
    pxcRom[4554] <= 10'b0000011100;
    pxcRom[4555] <= 10'b0000010000;
    pxcRom[4556] <= 10'b0000001001;
    pxcRom[4557] <= 10'b0000000100;
    pxcRom[4558] <= 10'b0000000001;
    pxcRom[4559] <= 10'b0000000000;
    pxcRom[4560] <= 10'b0000000000;
    pxcRom[4561] <= 10'b0000000000;
    pxcRom[4562] <= 10'b0000000000;
    pxcRom[4563] <= 10'b0000000000;
    pxcRom[4564] <= 10'b0000000000;
    pxcRom[4565] <= 10'b0000000000;
    pxcRom[4566] <= 10'b0000000000;
    pxcRom[4567] <= 10'b0000000000;
    pxcRom[4568] <= 10'b0000000000;
    pxcRom[4569] <= 10'b0000000010;
    pxcRom[4570] <= 10'b0000000111;
    pxcRom[4571] <= 10'b0000001111;
    pxcRom[4572] <= 10'b0000011010;
    pxcRom[4573] <= 10'b0000101000;
    pxcRom[4574] <= 10'b0000110110;
    pxcRom[4575] <= 10'b0001000001;
    pxcRom[4576] <= 10'b0001000011;
    pxcRom[4577] <= 10'b0001000001;
    pxcRom[4578] <= 10'b0000111011;
    pxcRom[4579] <= 10'b0000110000;
    pxcRom[4580] <= 10'b0000100100;
    pxcRom[4581] <= 10'b0000011000;
    pxcRom[4582] <= 10'b0000001110;
    pxcRom[4583] <= 10'b0000001000;
    pxcRom[4584] <= 10'b0000000100;
    pxcRom[4585] <= 10'b0000000001;
    pxcRom[4586] <= 10'b0000000000;
    pxcRom[4587] <= 10'b0000000000;
    pxcRom[4588] <= 10'b0000000000;
    pxcRom[4589] <= 10'b0000000000;
    pxcRom[4590] <= 10'b0000000000;
    pxcRom[4591] <= 10'b0000000000;
    pxcRom[4592] <= 10'b0000000000;
    pxcRom[4593] <= 10'b0000000000;
    pxcRom[4594] <= 10'b0000000000;
    pxcRom[4595] <= 10'b0000000000;
    pxcRom[4596] <= 10'b0000000000;
    pxcRom[4597] <= 10'b0000000000;
    pxcRom[4598] <= 10'b0000000010;
    pxcRom[4599] <= 10'b0000000101;
    pxcRom[4600] <= 10'b0000001001;
    pxcRom[4601] <= 10'b0000001111;
    pxcRom[4602] <= 10'b0000010101;
    pxcRom[4603] <= 10'b0000011001;
    pxcRom[4604] <= 10'b0000011100;
    pxcRom[4605] <= 10'b0000011011;
    pxcRom[4606] <= 10'b0000010111;
    pxcRom[4607] <= 10'b0000010010;
    pxcRom[4608] <= 10'b0000001100;
    pxcRom[4609] <= 10'b0000000111;
    pxcRom[4610] <= 10'b0000000100;
    pxcRom[4611] <= 10'b0000000010;
    pxcRom[4612] <= 10'b0000000001;
    pxcRom[4613] <= 10'b0000000000;
    pxcRom[4614] <= 10'b0000000000;
    pxcRom[4615] <= 10'b0000000000;
    pxcRom[4616] <= 10'b0000000000;
    pxcRom[4617] <= 10'b0000000000;
    pxcRom[4618] <= 10'b0000000000;
    pxcRom[4619] <= 10'b0000000000;
    pxcRom[4620] <= 10'b0000000000;
    pxcRom[4621] <= 10'b0000000000;
    pxcRom[4622] <= 10'b0000000000;
    pxcRom[4623] <= 10'b0000000000;
    pxcRom[4624] <= 10'b0000000000;
    pxcRom[4625] <= 10'b0000000000;
    pxcRom[4626] <= 10'b0000000000;
    pxcRom[4627] <= 10'b0000000000;
    pxcRom[4628] <= 10'b0000000001;
    pxcRom[4629] <= 10'b0000000010;
    pxcRom[4630] <= 10'b0000000011;
    pxcRom[4631] <= 10'b0000000100;
    pxcRom[4632] <= 10'b0000000100;
    pxcRom[4633] <= 10'b0000000100;
    pxcRom[4634] <= 10'b0000000011;
    pxcRom[4635] <= 10'b0000000010;
    pxcRom[4636] <= 10'b0000000001;
    pxcRom[4637] <= 10'b0000000001;
    pxcRom[4638] <= 10'b0000000000;
    pxcRom[4639] <= 10'b0000000000;
    pxcRom[4640] <= 10'b0000000000;
    pxcRom[4641] <= 10'b0000000000;
    pxcRom[4642] <= 10'b0000000000;
    pxcRom[4643] <= 10'b0000000000;
    pxcRom[4644] <= 10'b0000000000;
    pxcRom[4645] <= 10'b0000000000;
    pxcRom[4646] <= 10'b0000000000;
    pxcRom[4647] <= 10'b0000000000;
    pxcRom[4648] <= 10'b0000000000;
    pxcRom[4649] <= 10'b0000000000;
    pxcRom[4650] <= 10'b0000000000;
    pxcRom[4651] <= 10'b0000000000;
    pxcRom[4652] <= 10'b0000000000;
    pxcRom[4653] <= 10'b0000000000;
    pxcRom[4654] <= 10'b0000000000;
    pxcRom[4655] <= 10'b0000000000;
    pxcRom[4656] <= 10'b0000000000;
    pxcRom[4657] <= 10'b0000000000;
    pxcRom[4658] <= 10'b0000000000;
    pxcRom[4659] <= 10'b0000000000;
    pxcRom[4660] <= 10'b0000000000;
    pxcRom[4661] <= 10'b0000000000;
    pxcRom[4662] <= 10'b0000000000;
    pxcRom[4663] <= 10'b0000000000;
    pxcRom[4664] <= 10'b0000000000;
    pxcRom[4665] <= 10'b0000000000;
    pxcRom[4666] <= 10'b0000000000;
    pxcRom[4667] <= 10'b0000000000;
    pxcRom[4668] <= 10'b0000000000;
    pxcRom[4669] <= 10'b0000000000;
    pxcRom[4670] <= 10'b0000000000;
    pxcRom[4671] <= 10'b0000000000;
    pxcRom[4672] <= 10'b0000000000;
    pxcRom[4673] <= 10'b0000000000;
    pxcRom[4674] <= 10'b0000000000;
    pxcRom[4675] <= 10'b0000000000;
    pxcRom[4676] <= 10'b0000000000;
    pxcRom[4677] <= 10'b0000000000;
    pxcRom[4678] <= 10'b0000000000;
    pxcRom[4679] <= 10'b0000000000;
    pxcRom[4680] <= 10'b0000000000;
    pxcRom[4681] <= 10'b0000000000;
    pxcRom[4682] <= 10'b0000000000;
    pxcRom[4683] <= 10'b0000000000;
    pxcRom[4684] <= 10'b0000000000;
    pxcRom[4685] <= 10'b0000000000;
    pxcRom[4686] <= 10'b0000000000;
    pxcRom[4687] <= 10'b0000000000;
    pxcRom[4688] <= 10'b0000000000;
    pxcRom[4689] <= 10'b0000000000;
    pxcRom[4690] <= 10'b0000000000;
    pxcRom[4691] <= 10'b0000000000;
    pxcRom[4692] <= 10'b0000000000;
    pxcRom[4693] <= 10'b0000000000;
    pxcRom[4694] <= 10'b0000000000;
    pxcRom[4695] <= 10'b0000000000;
    pxcRom[4696] <= 10'b0000000000;
    pxcRom[4697] <= 10'b0000000000;
    pxcRom[4698] <= 10'b0000000000;
    pxcRom[4699] <= 10'b0000000000;
    pxcRom[4700] <= 10'b0000000000;
    pxcRom[4701] <= 10'b0000000000;
    pxcRom[4702] <= 10'b0000000000;
    pxcRom[4703] <= 10'b0000000000;
    pxcRom[4704] <= 10'b0000000000;
    pxcRom[4705] <= 10'b0000000000;
    pxcRom[4706] <= 10'b0000000000;
    pxcRom[4707] <= 10'b0000000000;
    pxcRom[4708] <= 10'b0000000000;
    pxcRom[4709] <= 10'b0000000000;
    pxcRom[4710] <= 10'b0000000000;
    pxcRom[4711] <= 10'b0000000000;
    pxcRom[4712] <= 10'b0000000000;
    pxcRom[4713] <= 10'b0000000000;
    pxcRom[4714] <= 10'b0000000000;
    pxcRom[4715] <= 10'b0000000000;
    pxcRom[4716] <= 10'b0000000000;
    pxcRom[4717] <= 10'b0000000000;
    pxcRom[4718] <= 10'b0000000000;
    pxcRom[4719] <= 10'b0000000000;
    pxcRom[4720] <= 10'b0000000000;
    pxcRom[4721] <= 10'b0000000000;
    pxcRom[4722] <= 10'b0000000000;
    pxcRom[4723] <= 10'b0000000000;
    pxcRom[4724] <= 10'b0000000000;
    pxcRom[4725] <= 10'b0000000000;
    pxcRom[4726] <= 10'b0000000000;
    pxcRom[4727] <= 10'b0000000000;
    pxcRom[4728] <= 10'b0000000000;
    pxcRom[4729] <= 10'b0000000000;
    pxcRom[4730] <= 10'b0000000000;
    pxcRom[4731] <= 10'b0000000000;
    pxcRom[4732] <= 10'b0000000000;
    pxcRom[4733] <= 10'b0000000000;
    pxcRom[4734] <= 10'b0000000000;
    pxcRom[4735] <= 10'b0000000000;
    pxcRom[4736] <= 10'b0000000000;
    pxcRom[4737] <= 10'b0000000000;
    pxcRom[4738] <= 10'b0000000000;
    pxcRom[4739] <= 10'b0000000000;
    pxcRom[4740] <= 10'b0000000000;
    pxcRom[4741] <= 10'b0000000000;
    pxcRom[4742] <= 10'b0000000000;
    pxcRom[4743] <= 10'b0000000000;
    pxcRom[4744] <= 10'b0000000000;
    pxcRom[4745] <= 10'b0000000000;
    pxcRom[4746] <= 10'b0000000000;
    pxcRom[4747] <= 10'b0000000000;
    pxcRom[4748] <= 10'b0000000000;
    pxcRom[4749] <= 10'b0000000000;
    pxcRom[4750] <= 10'b0000000000;
    pxcRom[4751] <= 10'b0000000000;
    pxcRom[4752] <= 10'b0000000000;
    pxcRom[4753] <= 10'b0000000000;
    pxcRom[4754] <= 10'b0000000000;
    pxcRom[4755] <= 10'b0000000000;
    pxcRom[4756] <= 10'b0000000000;
    pxcRom[4757] <= 10'b0000000000;
    pxcRom[4758] <= 10'b0000000000;
    pxcRom[4759] <= 10'b0000000000;
    pxcRom[4760] <= 10'b0000000000;
    pxcRom[4761] <= 10'b0000000000;
    pxcRom[4762] <= 10'b0000000000;
    pxcRom[4763] <= 10'b0000000000;
    pxcRom[4764] <= 10'b0000000000;
    pxcRom[4765] <= 10'b0000000000;
    pxcRom[4766] <= 10'b0000000000;
    pxcRom[4767] <= 10'b0000000000;
    pxcRom[4768] <= 10'b0000000000;
    pxcRom[4769] <= 10'b0000000001;
    pxcRom[4770] <= 10'b0000000010;
    pxcRom[4771] <= 10'b0000000100;
    pxcRom[4772] <= 10'b0000000110;
    pxcRom[4773] <= 10'b0000001000;
    pxcRom[4774] <= 10'b0000001011;
    pxcRom[4775] <= 10'b0000001101;
    pxcRom[4776] <= 10'b0000001110;
    pxcRom[4777] <= 10'b0000001100;
    pxcRom[4778] <= 10'b0000001010;
    pxcRom[4779] <= 10'b0000000111;
    pxcRom[4780] <= 10'b0000000100;
    pxcRom[4781] <= 10'b0000000010;
    pxcRom[4782] <= 10'b0000000001;
    pxcRom[4783] <= 10'b0000000000;
    pxcRom[4784] <= 10'b0000000000;
    pxcRom[4785] <= 10'b0000000000;
    pxcRom[4786] <= 10'b0000000000;
    pxcRom[4787] <= 10'b0000000000;
    pxcRom[4788] <= 10'b0000000000;
    pxcRom[4789] <= 10'b0000000000;
    pxcRom[4790] <= 10'b0000000000;
    pxcRom[4791] <= 10'b0000000000;
    pxcRom[4792] <= 10'b0000000000;
    pxcRom[4793] <= 10'b0000000000;
    pxcRom[4794] <= 10'b0000000000;
    pxcRom[4795] <= 10'b0000000000;
    pxcRom[4796] <= 10'b0000000001;
    pxcRom[4797] <= 10'b0000000011;
    pxcRom[4798] <= 10'b0000000101;
    pxcRom[4799] <= 10'b0000001000;
    pxcRom[4800] <= 10'b0000001101;
    pxcRom[4801] <= 10'b0000010011;
    pxcRom[4802] <= 10'b0000011011;
    pxcRom[4803] <= 10'b0000100001;
    pxcRom[4804] <= 10'b0000100101;
    pxcRom[4805] <= 10'b0000100011;
    pxcRom[4806] <= 10'b0000011101;
    pxcRom[4807] <= 10'b0000010100;
    pxcRom[4808] <= 10'b0000001011;
    pxcRom[4809] <= 10'b0000000101;
    pxcRom[4810] <= 10'b0000000011;
    pxcRom[4811] <= 10'b0000000001;
    pxcRom[4812] <= 10'b0000000000;
    pxcRom[4813] <= 10'b0000000000;
    pxcRom[4814] <= 10'b0000000000;
    pxcRom[4815] <= 10'b0000000000;
    pxcRom[4816] <= 10'b0000000000;
    pxcRom[4817] <= 10'b0000000000;
    pxcRom[4818] <= 10'b0000000000;
    pxcRom[4819] <= 10'b0000000000;
    pxcRom[4820] <= 10'b0000000000;
    pxcRom[4821] <= 10'b0000000000;
    pxcRom[4822] <= 10'b0000000000;
    pxcRom[4823] <= 10'b0000000001;
    pxcRom[4824] <= 10'b0000000010;
    pxcRom[4825] <= 10'b0000000100;
    pxcRom[4826] <= 10'b0000001000;
    pxcRom[4827] <= 10'b0000001100;
    pxcRom[4828] <= 10'b0000010100;
    pxcRom[4829] <= 10'b0000011100;
    pxcRom[4830] <= 10'b0000100111;
    pxcRom[4831] <= 10'b0000110000;
    pxcRom[4832] <= 10'b0000110011;
    pxcRom[4833] <= 10'b0000101100;
    pxcRom[4834] <= 10'b0000100001;
    pxcRom[4835] <= 10'b0000010110;
    pxcRom[4836] <= 10'b0000001100;
    pxcRom[4837] <= 10'b0000000110;
    pxcRom[4838] <= 10'b0000000011;
    pxcRom[4839] <= 10'b0000000001;
    pxcRom[4840] <= 10'b0000000000;
    pxcRom[4841] <= 10'b0000000000;
    pxcRom[4842] <= 10'b0000000000;
    pxcRom[4843] <= 10'b0000000000;
    pxcRom[4844] <= 10'b0000000000;
    pxcRom[4845] <= 10'b0000000000;
    pxcRom[4846] <= 10'b0000000000;
    pxcRom[4847] <= 10'b0000000000;
    pxcRom[4848] <= 10'b0000000000;
    pxcRom[4849] <= 10'b0000000000;
    pxcRom[4850] <= 10'b0000000000;
    pxcRom[4851] <= 10'b0000000001;
    pxcRom[4852] <= 10'b0000000011;
    pxcRom[4853] <= 10'b0000000111;
    pxcRom[4854] <= 10'b0000001011;
    pxcRom[4855] <= 10'b0000010010;
    pxcRom[4856] <= 10'b0000011100;
    pxcRom[4857] <= 10'b0000101000;
    pxcRom[4858] <= 10'b0000110010;
    pxcRom[4859] <= 10'b0000111001;
    pxcRom[4860] <= 10'b0000110011;
    pxcRom[4861] <= 10'b0000101000;
    pxcRom[4862] <= 10'b0000011011;
    pxcRom[4863] <= 10'b0000010000;
    pxcRom[4864] <= 10'b0000001001;
    pxcRom[4865] <= 10'b0000000100;
    pxcRom[4866] <= 10'b0000000010;
    pxcRom[4867] <= 10'b0000000001;
    pxcRom[4868] <= 10'b0000000000;
    pxcRom[4869] <= 10'b0000000000;
    pxcRom[4870] <= 10'b0000000000;
    pxcRom[4871] <= 10'b0000000000;
    pxcRom[4872] <= 10'b0000000000;
    pxcRom[4873] <= 10'b0000000000;
    pxcRom[4874] <= 10'b0000000000;
    pxcRom[4875] <= 10'b0000000000;
    pxcRom[4876] <= 10'b0000000000;
    pxcRom[4877] <= 10'b0000000000;
    pxcRom[4878] <= 10'b0000000001;
    pxcRom[4879] <= 10'b0000000010;
    pxcRom[4880] <= 10'b0000000101;
    pxcRom[4881] <= 10'b0000001001;
    pxcRom[4882] <= 10'b0000001111;
    pxcRom[4883] <= 10'b0000011001;
    pxcRom[4884] <= 10'b0000100101;
    pxcRom[4885] <= 10'b0000110011;
    pxcRom[4886] <= 10'b0000111011;
    pxcRom[4887] <= 10'b0000110111;
    pxcRom[4888] <= 10'b0000101010;
    pxcRom[4889] <= 10'b0000011100;
    pxcRom[4890] <= 10'b0000010001;
    pxcRom[4891] <= 10'b0000001001;
    pxcRom[4892] <= 10'b0000000101;
    pxcRom[4893] <= 10'b0000000010;
    pxcRom[4894] <= 10'b0000000001;
    pxcRom[4895] <= 10'b0000000000;
    pxcRom[4896] <= 10'b0000000000;
    pxcRom[4897] <= 10'b0000000000;
    pxcRom[4898] <= 10'b0000000000;
    pxcRom[4899] <= 10'b0000000000;
    pxcRom[4900] <= 10'b0000000000;
    pxcRom[4901] <= 10'b0000000000;
    pxcRom[4902] <= 10'b0000000000;
    pxcRom[4903] <= 10'b0000000000;
    pxcRom[4904] <= 10'b0000000000;
    pxcRom[4905] <= 10'b0000000000;
    pxcRom[4906] <= 10'b0000000001;
    pxcRom[4907] <= 10'b0000000011;
    pxcRom[4908] <= 10'b0000000111;
    pxcRom[4909] <= 10'b0000001100;
    pxcRom[4910] <= 10'b0000010101;
    pxcRom[4911] <= 10'b0000100010;
    pxcRom[4912] <= 10'b0000110000;
    pxcRom[4913] <= 10'b0000111100;
    pxcRom[4914] <= 10'b0000111011;
    pxcRom[4915] <= 10'b0000101110;
    pxcRom[4916] <= 10'b0000011101;
    pxcRom[4917] <= 10'b0000010001;
    pxcRom[4918] <= 10'b0000001001;
    pxcRom[4919] <= 10'b0000000100;
    pxcRom[4920] <= 10'b0000000010;
    pxcRom[4921] <= 10'b0000000001;
    pxcRom[4922] <= 10'b0000000000;
    pxcRom[4923] <= 10'b0000000000;
    pxcRom[4924] <= 10'b0000000000;
    pxcRom[4925] <= 10'b0000000000;
    pxcRom[4926] <= 10'b0000000000;
    pxcRom[4927] <= 10'b0000000000;
    pxcRom[4928] <= 10'b0000000000;
    pxcRom[4929] <= 10'b0000000000;
    pxcRom[4930] <= 10'b0000000000;
    pxcRom[4931] <= 10'b0000000000;
    pxcRom[4932] <= 10'b0000000000;
    pxcRom[4933] <= 10'b0000000000;
    pxcRom[4934] <= 10'b0000000001;
    pxcRom[4935] <= 10'b0000000100;
    pxcRom[4936] <= 10'b0000001001;
    pxcRom[4937] <= 10'b0000010001;
    pxcRom[4938] <= 10'b0000011101;
    pxcRom[4939] <= 10'b0000101100;
    pxcRom[4940] <= 10'b0000111100;
    pxcRom[4941] <= 10'b0001000001;
    pxcRom[4942] <= 10'b0000110100;
    pxcRom[4943] <= 10'b0000100010;
    pxcRom[4944] <= 10'b0000010010;
    pxcRom[4945] <= 10'b0000001001;
    pxcRom[4946] <= 10'b0000000100;
    pxcRom[4947] <= 10'b0000000010;
    pxcRom[4948] <= 10'b0000000010;
    pxcRom[4949] <= 10'b0000000001;
    pxcRom[4950] <= 10'b0000000000;
    pxcRom[4951] <= 10'b0000000000;
    pxcRom[4952] <= 10'b0000000000;
    pxcRom[4953] <= 10'b0000000000;
    pxcRom[4954] <= 10'b0000000000;
    pxcRom[4955] <= 10'b0000000000;
    pxcRom[4956] <= 10'b0000000000;
    pxcRom[4957] <= 10'b0000000000;
    pxcRom[4958] <= 10'b0000000000;
    pxcRom[4959] <= 10'b0000000000;
    pxcRom[4960] <= 10'b0000000000;
    pxcRom[4961] <= 10'b0000000000;
    pxcRom[4962] <= 10'b0000000010;
    pxcRom[4963] <= 10'b0000000110;
    pxcRom[4964] <= 10'b0000001100;
    pxcRom[4965] <= 10'b0000010111;
    pxcRom[4966] <= 10'b0000100110;
    pxcRom[4967] <= 10'b0000111001;
    pxcRom[4968] <= 10'b0001000101;
    pxcRom[4969] <= 10'b0000111101;
    pxcRom[4970] <= 10'b0000101001;
    pxcRom[4971] <= 10'b0000010110;
    pxcRom[4972] <= 10'b0000001011;
    pxcRom[4973] <= 10'b0000000101;
    pxcRom[4974] <= 10'b0000000011;
    pxcRom[4975] <= 10'b0000000011;
    pxcRom[4976] <= 10'b0000000011;
    pxcRom[4977] <= 10'b0000000010;
    pxcRom[4978] <= 10'b0000000001;
    pxcRom[4979] <= 10'b0000000000;
    pxcRom[4980] <= 10'b0000000000;
    pxcRom[4981] <= 10'b0000000000;
    pxcRom[4982] <= 10'b0000000000;
    pxcRom[4983] <= 10'b0000000000;
    pxcRom[4984] <= 10'b0000000000;
    pxcRom[4985] <= 10'b0000000000;
    pxcRom[4986] <= 10'b0000000000;
    pxcRom[4987] <= 10'b0000000000;
    pxcRom[4988] <= 10'b0000000000;
    pxcRom[4989] <= 10'b0000000000;
    pxcRom[4990] <= 10'b0000000011;
    pxcRom[4991] <= 10'b0000001000;
    pxcRom[4992] <= 10'b0000010000;
    pxcRom[4993] <= 10'b0000011111;
    pxcRom[4994] <= 10'b0000110010;
    pxcRom[4995] <= 10'b0001000110;
    pxcRom[4996] <= 10'b0001000111;
    pxcRom[4997] <= 10'b0000110100;
    pxcRom[4998] <= 10'b0000011101;
    pxcRom[4999] <= 10'b0000001111;
    pxcRom[5000] <= 10'b0000001001;
    pxcRom[5001] <= 10'b0000000111;
    pxcRom[5002] <= 10'b0000001000;
    pxcRom[5003] <= 10'b0000001000;
    pxcRom[5004] <= 10'b0000001000;
    pxcRom[5005] <= 10'b0000000110;
    pxcRom[5006] <= 10'b0000000100;
    pxcRom[5007] <= 10'b0000000001;
    pxcRom[5008] <= 10'b0000000000;
    pxcRom[5009] <= 10'b0000000000;
    pxcRom[5010] <= 10'b0000000000;
    pxcRom[5011] <= 10'b0000000000;
    pxcRom[5012] <= 10'b0000000000;
    pxcRom[5013] <= 10'b0000000000;
    pxcRom[5014] <= 10'b0000000000;
    pxcRom[5015] <= 10'b0000000000;
    pxcRom[5016] <= 10'b0000000000;
    pxcRom[5017] <= 10'b0000000001;
    pxcRom[5018] <= 10'b0000000100;
    pxcRom[5019] <= 10'b0000001010;
    pxcRom[5020] <= 10'b0000010110;
    pxcRom[5021] <= 10'b0000101001;
    pxcRom[5022] <= 10'b0001000000;
    pxcRom[5023] <= 10'b0001001110;
    pxcRom[5024] <= 10'b0001000011;
    pxcRom[5025] <= 10'b0000101010;
    pxcRom[5026] <= 10'b0000010111;
    pxcRom[5027] <= 10'b0000001110;
    pxcRom[5028] <= 10'b0000001111;
    pxcRom[5029] <= 10'b0000010010;
    pxcRom[5030] <= 10'b0000010100;
    pxcRom[5031] <= 10'b0000010100;
    pxcRom[5032] <= 10'b0000010001;
    pxcRom[5033] <= 10'b0000001100;
    pxcRom[5034] <= 10'b0000000111;
    pxcRom[5035] <= 10'b0000000100;
    pxcRom[5036] <= 10'b0000000001;
    pxcRom[5037] <= 10'b0000000000;
    pxcRom[5038] <= 10'b0000000000;
    pxcRom[5039] <= 10'b0000000000;
    pxcRom[5040] <= 10'b0000000000;
    pxcRom[5041] <= 10'b0000000000;
    pxcRom[5042] <= 10'b0000000000;
    pxcRom[5043] <= 10'b0000000000;
    pxcRom[5044] <= 10'b0000000000;
    pxcRom[5045] <= 10'b0000000001;
    pxcRom[5046] <= 10'b0000000101;
    pxcRom[5047] <= 10'b0000001101;
    pxcRom[5048] <= 10'b0000011100;
    pxcRom[5049] <= 10'b0000110101;
    pxcRom[5050] <= 10'b0001010000;
    pxcRom[5051] <= 10'b0001010001;
    pxcRom[5052] <= 10'b0000111001;
    pxcRom[5053] <= 10'b0000100011;
    pxcRom[5054] <= 10'b0000011000;
    pxcRom[5055] <= 10'b0000011010;
    pxcRom[5056] <= 10'b0000100010;
    pxcRom[5057] <= 10'b0000101000;
    pxcRom[5058] <= 10'b0000101001;
    pxcRom[5059] <= 10'b0000100110;
    pxcRom[5060] <= 10'b0000011111;
    pxcRom[5061] <= 10'b0000010110;
    pxcRom[5062] <= 10'b0000001110;
    pxcRom[5063] <= 10'b0000000111;
    pxcRom[5064] <= 10'b0000000011;
    pxcRom[5065] <= 10'b0000000000;
    pxcRom[5066] <= 10'b0000000000;
    pxcRom[5067] <= 10'b0000000000;
    pxcRom[5068] <= 10'b0000000000;
    pxcRom[5069] <= 10'b0000000000;
    pxcRom[5070] <= 10'b0000000000;
    pxcRom[5071] <= 10'b0000000000;
    pxcRom[5072] <= 10'b0000000000;
    pxcRom[5073] <= 10'b0000000001;
    pxcRom[5074] <= 10'b0000000111;
    pxcRom[5075] <= 10'b0000010001;
    pxcRom[5076] <= 10'b0000100101;
    pxcRom[5077] <= 10'b0001000001;
    pxcRom[5078] <= 10'b0001011001;
    pxcRom[5079] <= 10'b0001001110;
    pxcRom[5080] <= 10'b0000110011;
    pxcRom[5081] <= 10'b0000100101;
    pxcRom[5082] <= 10'b0000100111;
    pxcRom[5083] <= 10'b0000110100;
    pxcRom[5084] <= 10'b0001000010;
    pxcRom[5085] <= 10'b0001000111;
    pxcRom[5086] <= 10'b0001000010;
    pxcRom[5087] <= 10'b0000111010;
    pxcRom[5088] <= 10'b0000101101;
    pxcRom[5089] <= 10'b0000100000;
    pxcRom[5090] <= 10'b0000010100;
    pxcRom[5091] <= 10'b0000001010;
    pxcRom[5092] <= 10'b0000000100;
    pxcRom[5093] <= 10'b0000000000;
    pxcRom[5094] <= 10'b0000000000;
    pxcRom[5095] <= 10'b0000000000;
    pxcRom[5096] <= 10'b0000000000;
    pxcRom[5097] <= 10'b0000000000;
    pxcRom[5098] <= 10'b0000000000;
    pxcRom[5099] <= 10'b0000000000;
    pxcRom[5100] <= 10'b0000000000;
    pxcRom[5101] <= 10'b0000000010;
    pxcRom[5102] <= 10'b0000001000;
    pxcRom[5103] <= 10'b0000010110;
    pxcRom[5104] <= 10'b0000101101;
    pxcRom[5105] <= 10'b0001010000;
    pxcRom[5106] <= 10'b0001100000;
    pxcRom[5107] <= 10'b0001001001;
    pxcRom[5108] <= 10'b0000110011;
    pxcRom[5109] <= 10'b0000110000;
    pxcRom[5110] <= 10'b0000111111;
    pxcRom[5111] <= 10'b0001010100;
    pxcRom[5112] <= 10'b0001011101;
    pxcRom[5113] <= 10'b0001010111;
    pxcRom[5114] <= 10'b0001001011;
    pxcRom[5115] <= 10'b0001000100;
    pxcRom[5116] <= 10'b0000111000;
    pxcRom[5117] <= 10'b0000101001;
    pxcRom[5118] <= 10'b0000011001;
    pxcRom[5119] <= 10'b0000001101;
    pxcRom[5120] <= 10'b0000000101;
    pxcRom[5121] <= 10'b0000000001;
    pxcRom[5122] <= 10'b0000000000;
    pxcRom[5123] <= 10'b0000000000;
    pxcRom[5124] <= 10'b0000000000;
    pxcRom[5125] <= 10'b0000000000;
    pxcRom[5126] <= 10'b0000000000;
    pxcRom[5127] <= 10'b0000000000;
    pxcRom[5128] <= 10'b0000000000;
    pxcRom[5129] <= 10'b0000000010;
    pxcRom[5130] <= 10'b0000001010;
    pxcRom[5131] <= 10'b0000011010;
    pxcRom[5132] <= 10'b0000110101;
    pxcRom[5133] <= 10'b0001011001;
    pxcRom[5134] <= 10'b0001100010;
    pxcRom[5135] <= 10'b0001001000;
    pxcRom[5136] <= 10'b0000111000;
    pxcRom[5137] <= 10'b0001000000;
    pxcRom[5138] <= 10'b0001010100;
    pxcRom[5139] <= 10'b0001011011;
    pxcRom[5140] <= 10'b0001001111;
    pxcRom[5141] <= 10'b0001000100;
    pxcRom[5142] <= 10'b0001000001;
    pxcRom[5143] <= 10'b0001000011;
    pxcRom[5144] <= 10'b0000111110;
    pxcRom[5145] <= 10'b0000101110;
    pxcRom[5146] <= 10'b0000011100;
    pxcRom[5147] <= 10'b0000001110;
    pxcRom[5148] <= 10'b0000000110;
    pxcRom[5149] <= 10'b0000000001;
    pxcRom[5150] <= 10'b0000000000;
    pxcRom[5151] <= 10'b0000000000;
    pxcRom[5152] <= 10'b0000000000;
    pxcRom[5153] <= 10'b0000000000;
    pxcRom[5154] <= 10'b0000000000;
    pxcRom[5155] <= 10'b0000000000;
    pxcRom[5156] <= 10'b0000000000;
    pxcRom[5157] <= 10'b0000000011;
    pxcRom[5158] <= 10'b0000001011;
    pxcRom[5159] <= 10'b0000011100;
    pxcRom[5160] <= 10'b0000111011;
    pxcRom[5161] <= 10'b0001011111;
    pxcRom[5162] <= 10'b0001100101;
    pxcRom[5163] <= 10'b0001001101;
    pxcRom[5164] <= 10'b0001000010;
    pxcRom[5165] <= 10'b0001001000;
    pxcRom[5166] <= 10'b0001001110;
    pxcRom[5167] <= 10'b0001000010;
    pxcRom[5168] <= 10'b0000110100;
    pxcRom[5169] <= 10'b0000110001;
    pxcRom[5170] <= 10'b0000111011;
    pxcRom[5171] <= 10'b0001001001;
    pxcRom[5172] <= 10'b0001000100;
    pxcRom[5173] <= 10'b0000101111;
    pxcRom[5174] <= 10'b0000011011;
    pxcRom[5175] <= 10'b0000001100;
    pxcRom[5176] <= 10'b0000000101;
    pxcRom[5177] <= 10'b0000000001;
    pxcRom[5178] <= 10'b0000000000;
    pxcRom[5179] <= 10'b0000000000;
    pxcRom[5180] <= 10'b0000000000;
    pxcRom[5181] <= 10'b0000000000;
    pxcRom[5182] <= 10'b0000000000;
    pxcRom[5183] <= 10'b0000000000;
    pxcRom[5184] <= 10'b0000000000;
    pxcRom[5185] <= 10'b0000000011;
    pxcRom[5186] <= 10'b0000001011;
    pxcRom[5187] <= 10'b0000011100;
    pxcRom[5188] <= 10'b0000111011;
    pxcRom[5189] <= 10'b0001100000;
    pxcRom[5190] <= 10'b0001110000;
    pxcRom[5191] <= 10'b0001011011;
    pxcRom[5192] <= 10'b0001001010;
    pxcRom[5193] <= 10'b0001000110;
    pxcRom[5194] <= 10'b0000111101;
    pxcRom[5195] <= 10'b0000110000;
    pxcRom[5196] <= 10'b0000101100;
    pxcRom[5197] <= 10'b0000110101;
    pxcRom[5198] <= 10'b0001001000;
    pxcRom[5199] <= 10'b0001010101;
    pxcRom[5200] <= 10'b0001000101;
    pxcRom[5201] <= 10'b0000101011;
    pxcRom[5202] <= 10'b0000010110;
    pxcRom[5203] <= 10'b0000001001;
    pxcRom[5204] <= 10'b0000000100;
    pxcRom[5205] <= 10'b0000000001;
    pxcRom[5206] <= 10'b0000000000;
    pxcRom[5207] <= 10'b0000000000;
    pxcRom[5208] <= 10'b0000000000;
    pxcRom[5209] <= 10'b0000000000;
    pxcRom[5210] <= 10'b0000000000;
    pxcRom[5211] <= 10'b0000000000;
    pxcRom[5212] <= 10'b0000000000;
    pxcRom[5213] <= 10'b0000000010;
    pxcRom[5214] <= 10'b0000001001;
    pxcRom[5215] <= 10'b0000011001;
    pxcRom[5216] <= 10'b0000110101;
    pxcRom[5217] <= 10'b0001100000;
    pxcRom[5218] <= 10'b0010000001;
    pxcRom[5219] <= 10'b0001110100;
    pxcRom[5220] <= 10'b0001011000;
    pxcRom[5221] <= 10'b0001000111;
    pxcRom[5222] <= 10'b0000111100;
    pxcRom[5223] <= 10'b0000111010;
    pxcRom[5224] <= 10'b0001000001;
    pxcRom[5225] <= 10'b0001010101;
    pxcRom[5226] <= 10'b0001100111;
    pxcRom[5227] <= 10'b0001011001;
    pxcRom[5228] <= 10'b0000111010;
    pxcRom[5229] <= 10'b0000100000;
    pxcRom[5230] <= 10'b0000001111;
    pxcRom[5231] <= 10'b0000000110;
    pxcRom[5232] <= 10'b0000000010;
    pxcRom[5233] <= 10'b0000000000;
    pxcRom[5234] <= 10'b0000000000;
    pxcRom[5235] <= 10'b0000000000;
    pxcRom[5236] <= 10'b0000000000;
    pxcRom[5237] <= 10'b0000000000;
    pxcRom[5238] <= 10'b0000000000;
    pxcRom[5239] <= 10'b0000000000;
    pxcRom[5240] <= 10'b0000000000;
    pxcRom[5241] <= 10'b0000000001;
    pxcRom[5242] <= 10'b0000000110;
    pxcRom[5243] <= 10'b0000010011;
    pxcRom[5244] <= 10'b0000101010;
    pxcRom[5245] <= 10'b0001010010;
    pxcRom[5246] <= 10'b0010000101;
    pxcRom[5247] <= 10'b0010010111;
    pxcRom[5248] <= 10'b0001111100;
    pxcRom[5249] <= 10'b0001100101;
    pxcRom[5250] <= 10'b0001011101;
    pxcRom[5251] <= 10'b0001100100;
    pxcRom[5252] <= 10'b0001110011;
    pxcRom[5253] <= 10'b0001111111;
    pxcRom[5254] <= 10'b0001101010;
    pxcRom[5255] <= 10'b0001000100;
    pxcRom[5256] <= 10'b0000100111;
    pxcRom[5257] <= 10'b0000010011;
    pxcRom[5258] <= 10'b0000001001;
    pxcRom[5259] <= 10'b0000000011;
    pxcRom[5260] <= 10'b0000000001;
    pxcRom[5261] <= 10'b0000000000;
    pxcRom[5262] <= 10'b0000000000;
    pxcRom[5263] <= 10'b0000000000;
    pxcRom[5264] <= 10'b0000000000;
    pxcRom[5265] <= 10'b0000000000;
    pxcRom[5266] <= 10'b0000000000;
    pxcRom[5267] <= 10'b0000000000;
    pxcRom[5268] <= 10'b0000000000;
    pxcRom[5269] <= 10'b0000000001;
    pxcRom[5270] <= 10'b0000000011;
    pxcRom[5271] <= 10'b0000001011;
    pxcRom[5272] <= 10'b0000011011;
    pxcRom[5273] <= 10'b0000110111;
    pxcRom[5274] <= 10'b0001100101;
    pxcRom[5275] <= 10'b0010011001;
    pxcRom[5276] <= 10'b0010110101;
    pxcRom[5277] <= 10'b0010101001;
    pxcRom[5278] <= 10'b0010100100;
    pxcRom[5279] <= 10'b0010011111;
    pxcRom[5280] <= 10'b0010001010;
    pxcRom[5281] <= 10'b0001101001;
    pxcRom[5282] <= 10'b0001000011;
    pxcRom[5283] <= 10'b0000100110;
    pxcRom[5284] <= 10'b0000010011;
    pxcRom[5285] <= 10'b0000001001;
    pxcRom[5286] <= 10'b0000000011;
    pxcRom[5287] <= 10'b0000000001;
    pxcRom[5288] <= 10'b0000000000;
    pxcRom[5289] <= 10'b0000000000;
    pxcRom[5290] <= 10'b0000000000;
    pxcRom[5291] <= 10'b0000000000;
    pxcRom[5292] <= 10'b0000000000;
    pxcRom[5293] <= 10'b0000000000;
    pxcRom[5294] <= 10'b0000000000;
    pxcRom[5295] <= 10'b0000000000;
    pxcRom[5296] <= 10'b0000000000;
    pxcRom[5297] <= 10'b0000000000;
    pxcRom[5298] <= 10'b0000000001;
    pxcRom[5299] <= 10'b0000000101;
    pxcRom[5300] <= 10'b0000001100;
    pxcRom[5301] <= 10'b0000011100;
    pxcRom[5302] <= 10'b0000110100;
    pxcRom[5303] <= 10'b0001010110;
    pxcRom[5304] <= 10'b0001111000;
    pxcRom[5305] <= 10'b0010001000;
    pxcRom[5306] <= 10'b0001111111;
    pxcRom[5307] <= 10'b0001101000;
    pxcRom[5308] <= 10'b0001001100;
    pxcRom[5309] <= 10'b0000110001;
    pxcRom[5310] <= 10'b0000011101;
    pxcRom[5311] <= 10'b0000001111;
    pxcRom[5312] <= 10'b0000000111;
    pxcRom[5313] <= 10'b0000000010;
    pxcRom[5314] <= 10'b0000000001;
    pxcRom[5315] <= 10'b0000000000;
    pxcRom[5316] <= 10'b0000000000;
    pxcRom[5317] <= 10'b0000000000;
    pxcRom[5318] <= 10'b0000000000;
    pxcRom[5319] <= 10'b0000000000;
    pxcRom[5320] <= 10'b0000000000;
    pxcRom[5321] <= 10'b0000000000;
    pxcRom[5322] <= 10'b0000000000;
    pxcRom[5323] <= 10'b0000000000;
    pxcRom[5324] <= 10'b0000000000;
    pxcRom[5325] <= 10'b0000000000;
    pxcRom[5326] <= 10'b0000000000;
    pxcRom[5327] <= 10'b0000000001;
    pxcRom[5328] <= 10'b0000000011;
    pxcRom[5329] <= 10'b0000000110;
    pxcRom[5330] <= 10'b0000001100;
    pxcRom[5331] <= 10'b0000010100;
    pxcRom[5332] <= 10'b0000011011;
    pxcRom[5333] <= 10'b0000011110;
    pxcRom[5334] <= 10'b0000011101;
    pxcRom[5335] <= 10'b0000011000;
    pxcRom[5336] <= 10'b0000010010;
    pxcRom[5337] <= 10'b0000001011;
    pxcRom[5338] <= 10'b0000000110;
    pxcRom[5339] <= 10'b0000000011;
    pxcRom[5340] <= 10'b0000000001;
    pxcRom[5341] <= 10'b0000000000;
    pxcRom[5342] <= 10'b0000000000;
    pxcRom[5343] <= 10'b0000000000;
    pxcRom[5344] <= 10'b0000000000;
    pxcRom[5345] <= 10'b0000000000;
    pxcRom[5346] <= 10'b0000000000;
    pxcRom[5347] <= 10'b0000000000;
    pxcRom[5348] <= 10'b0000000000;
    pxcRom[5349] <= 10'b0000000000;
    pxcRom[5350] <= 10'b0000000000;
    pxcRom[5351] <= 10'b0000000000;
    pxcRom[5352] <= 10'b0000000000;
    pxcRom[5353] <= 10'b0000000000;
    pxcRom[5354] <= 10'b0000000000;
    pxcRom[5355] <= 10'b0000000000;
    pxcRom[5356] <= 10'b0000000000;
    pxcRom[5357] <= 10'b0000000000;
    pxcRom[5358] <= 10'b0000000000;
    pxcRom[5359] <= 10'b0000000001;
    pxcRom[5360] <= 10'b0000000010;
    pxcRom[5361] <= 10'b0000000010;
    pxcRom[5362] <= 10'b0000000010;
    pxcRom[5363] <= 10'b0000000010;
    pxcRom[5364] <= 10'b0000000001;
    pxcRom[5365] <= 10'b0000000001;
    pxcRom[5366] <= 10'b0000000000;
    pxcRom[5367] <= 10'b0000000000;
    pxcRom[5368] <= 10'b0000000000;
    pxcRom[5369] <= 10'b0000000000;
    pxcRom[5370] <= 10'b0000000000;
    pxcRom[5371] <= 10'b0000000000;
    pxcRom[5372] <= 10'b0000000000;
    pxcRom[5373] <= 10'b0000000000;
    pxcRom[5374] <= 10'b0000000000;
    pxcRom[5375] <= 10'b0000000000;
    pxcRom[5376] <= 10'b0000000000;
    pxcRom[5377] <= 10'b0000000000;
    pxcRom[5378] <= 10'b0000000000;
    pxcRom[5379] <= 10'b0000000000;
    pxcRom[5380] <= 10'b0000000000;
    pxcRom[5381] <= 10'b0000000000;
    pxcRom[5382] <= 10'b0000000000;
    pxcRom[5383] <= 10'b0000000000;
    pxcRom[5384] <= 10'b0000000000;
    pxcRom[5385] <= 10'b0000000000;
    pxcRom[5386] <= 10'b0000000000;
    pxcRom[5387] <= 10'b0000000000;
    pxcRom[5388] <= 10'b0000000000;
    pxcRom[5389] <= 10'b0000000000;
    pxcRom[5390] <= 10'b0000000000;
    pxcRom[5391] <= 10'b0000000000;
    pxcRom[5392] <= 10'b0000000000;
    pxcRom[5393] <= 10'b0000000000;
    pxcRom[5394] <= 10'b0000000000;
    pxcRom[5395] <= 10'b0000000000;
    pxcRom[5396] <= 10'b0000000000;
    pxcRom[5397] <= 10'b0000000000;
    pxcRom[5398] <= 10'b0000000000;
    pxcRom[5399] <= 10'b0000000000;
    pxcRom[5400] <= 10'b0000000000;
    pxcRom[5401] <= 10'b0000000000;
    pxcRom[5402] <= 10'b0000000000;
    pxcRom[5403] <= 10'b0000000000;
    pxcRom[5404] <= 10'b0000000000;
    pxcRom[5405] <= 10'b0000000000;
    pxcRom[5406] <= 10'b0000000000;
    pxcRom[5407] <= 10'b0000000000;
    pxcRom[5408] <= 10'b0000000000;
    pxcRom[5409] <= 10'b0000000000;
    pxcRom[5410] <= 10'b0000000000;
    pxcRom[5411] <= 10'b0000000000;
    pxcRom[5412] <= 10'b0000000000;
    pxcRom[5413] <= 10'b0000000000;
    pxcRom[5414] <= 10'b0000000000;
    pxcRom[5415] <= 10'b0000000000;
    pxcRom[5416] <= 10'b0000000000;
    pxcRom[5417] <= 10'b0000000000;
    pxcRom[5418] <= 10'b0000000000;
    pxcRom[5419] <= 10'b0000000000;
    pxcRom[5420] <= 10'b0000000000;
    pxcRom[5421] <= 10'b0000000000;
    pxcRom[5422] <= 10'b0000000000;
    pxcRom[5423] <= 10'b0000000000;
    pxcRom[5424] <= 10'b0000000000;
    pxcRom[5425] <= 10'b0000000000;
    pxcRom[5426] <= 10'b0000000000;
    pxcRom[5427] <= 10'b0000000000;
    pxcRom[5428] <= 10'b0000000000;
    pxcRom[5429] <= 10'b0000000000;
    pxcRom[5430] <= 10'b0000000000;
    pxcRom[5431] <= 10'b0000000000;
    pxcRom[5432] <= 10'b0000000000;
    pxcRom[5433] <= 10'b0000000000;
    pxcRom[5434] <= 10'b0000000000;
    pxcRom[5435] <= 10'b0000000000;
    pxcRom[5436] <= 10'b0000000000;
    pxcRom[5437] <= 10'b0000000000;
    pxcRom[5438] <= 10'b0000000000;
    pxcRom[5439] <= 10'b0000000000;
    pxcRom[5440] <= 10'b0000000000;
    pxcRom[5441] <= 10'b0000000000;
    pxcRom[5442] <= 10'b0000000000;
    pxcRom[5443] <= 10'b0000000000;
    pxcRom[5444] <= 10'b0000000000;
    pxcRom[5445] <= 10'b0000000000;
    pxcRom[5446] <= 10'b0000000000;
    pxcRom[5447] <= 10'b0000000000;
    pxcRom[5448] <= 10'b0000000000;
    pxcRom[5449] <= 10'b0000000000;
    pxcRom[5450] <= 10'b0000000000;
    pxcRom[5451] <= 10'b0000000000;
    pxcRom[5452] <= 10'b0000000000;
    pxcRom[5453] <= 10'b0000000000;
    pxcRom[5454] <= 10'b0000000000;
    pxcRom[5455] <= 10'b0000000000;
    pxcRom[5456] <= 10'b0000000000;
    pxcRom[5457] <= 10'b0000000000;
    pxcRom[5458] <= 10'b0000000000;
    pxcRom[5459] <= 10'b0000000000;
    pxcRom[5460] <= 10'b0000000000;
    pxcRom[5461] <= 10'b0000000000;
    pxcRom[5462] <= 10'b0000000000;
    pxcRom[5463] <= 10'b0000000000;
    pxcRom[5464] <= 10'b0000000000;
    pxcRom[5465] <= 10'b0000000000;
    pxcRom[5466] <= 10'b0000000000;
    pxcRom[5467] <= 10'b0000000000;
    pxcRom[5468] <= 10'b0000000000;
    pxcRom[5469] <= 10'b0000000000;
    pxcRom[5470] <= 10'b0000000000;
    pxcRom[5471] <= 10'b0000000000;
    pxcRom[5472] <= 10'b0000000000;
    pxcRom[5473] <= 10'b0000000000;
    pxcRom[5474] <= 10'b0000000000;
    pxcRom[5475] <= 10'b0000000000;
    pxcRom[5476] <= 10'b0000000000;
    pxcRom[5477] <= 10'b0000000000;
    pxcRom[5478] <= 10'b0000000000;
    pxcRom[5479] <= 10'b0000000000;
    pxcRom[5480] <= 10'b0000000000;
    pxcRom[5481] <= 10'b0000000000;
    pxcRom[5482] <= 10'b0000000000;
    pxcRom[5483] <= 10'b0000000000;
    pxcRom[5484] <= 10'b0000000000;
    pxcRom[5485] <= 10'b0000000000;
    pxcRom[5486] <= 10'b0000000000;
    pxcRom[5487] <= 10'b0000000000;
    pxcRom[5488] <= 10'b0000000000;
    pxcRom[5489] <= 10'b0000000000;
    pxcRom[5490] <= 10'b0000000000;
    pxcRom[5491] <= 10'b0000000000;
    pxcRom[5492] <= 10'b0000000000;
    pxcRom[5493] <= 10'b0000000000;
    pxcRom[5494] <= 10'b0000000000;
    pxcRom[5495] <= 10'b0000000000;
    pxcRom[5496] <= 10'b0000000000;
    pxcRom[5497] <= 10'b0000000000;
    pxcRom[5498] <= 10'b0000000000;
    pxcRom[5499] <= 10'b0000000000;
    pxcRom[5500] <= 10'b0000000000;
    pxcRom[5501] <= 10'b0000000000;
    pxcRom[5502] <= 10'b0000000000;
    pxcRom[5503] <= 10'b0000000000;
    pxcRom[5504] <= 10'b0000000000;
    pxcRom[5505] <= 10'b0000000000;
    pxcRom[5506] <= 10'b0000000000;
    pxcRom[5507] <= 10'b0000000000;
    pxcRom[5508] <= 10'b0000000000;
    pxcRom[5509] <= 10'b0000000000;
    pxcRom[5510] <= 10'b0000000000;
    pxcRom[5511] <= 10'b0000000000;
    pxcRom[5512] <= 10'b0000000000;
    pxcRom[5513] <= 10'b0000000000;
    pxcRom[5514] <= 10'b0000000000;
    pxcRom[5515] <= 10'b0000000000;
    pxcRom[5516] <= 10'b0000000000;
    pxcRom[5517] <= 10'b0000000000;
    pxcRom[5518] <= 10'b0000000000;
    pxcRom[5519] <= 10'b0000000000;
    pxcRom[5520] <= 10'b0000000000;
    pxcRom[5521] <= 10'b0000000000;
    pxcRom[5522] <= 10'b0000000000;
    pxcRom[5523] <= 10'b0000000000;
    pxcRom[5524] <= 10'b0000000000;
    pxcRom[5525] <= 10'b0000000000;
    pxcRom[5526] <= 10'b0000000000;
    pxcRom[5527] <= 10'b0000000000;
    pxcRom[5528] <= 10'b0000000000;
    pxcRom[5529] <= 10'b0000000000;
    pxcRom[5530] <= 10'b0000000000;
    pxcRom[5531] <= 10'b0000000000;
    pxcRom[5532] <= 10'b0000000000;
    pxcRom[5533] <= 10'b0000000000;
    pxcRom[5534] <= 10'b0000000000;
    pxcRom[5535] <= 10'b0000000000;
    pxcRom[5536] <= 10'b0000000000;
    pxcRom[5537] <= 10'b0000000000;
    pxcRom[5538] <= 10'b0000000000;
    pxcRom[5539] <= 10'b0000000000;
    pxcRom[5540] <= 10'b0000000000;
    pxcRom[5541] <= 10'b0000000000;
    pxcRom[5542] <= 10'b0000000000;
    pxcRom[5543] <= 10'b0000000000;
    pxcRom[5544] <= 10'b0000000000;
    pxcRom[5545] <= 10'b0000000000;
    pxcRom[5546] <= 10'b0000000000;
    pxcRom[5547] <= 10'b0000000000;
    pxcRom[5548] <= 10'b0000000000;
    pxcRom[5549] <= 10'b0000000000;
    pxcRom[5550] <= 10'b0000000000;
    pxcRom[5551] <= 10'b0000000000;
    pxcRom[5552] <= 10'b0000000000;
    pxcRom[5553] <= 10'b0000000000;
    pxcRom[5554] <= 10'b0000000000;
    pxcRom[5555] <= 10'b0000000000;
    pxcRom[5556] <= 10'b0000000000;
    pxcRom[5557] <= 10'b0000000000;
    pxcRom[5558] <= 10'b0000000000;
    pxcRom[5559] <= 10'b0000000000;
    pxcRom[5560] <= 10'b0000000000;
    pxcRom[5561] <= 10'b0000000000;
    pxcRom[5562] <= 10'b0000000000;
    pxcRom[5563] <= 10'b0000000000;
    pxcRom[5564] <= 10'b0000000000;
    pxcRom[5565] <= 10'b0000000000;
    pxcRom[5566] <= 10'b0000000000;
    pxcRom[5567] <= 10'b0000000000;
    pxcRom[5568] <= 10'b0000000000;
    pxcRom[5569] <= 10'b0000000000;
    pxcRom[5570] <= 10'b0000000000;
    pxcRom[5571] <= 10'b0000000000;
    pxcRom[5572] <= 10'b0000000000;
    pxcRom[5573] <= 10'b0000000000;
    pxcRom[5574] <= 10'b0000000000;
    pxcRom[5575] <= 10'b0000000000;
    pxcRom[5576] <= 10'b0000000000;
    pxcRom[5577] <= 10'b0000000000;
    pxcRom[5578] <= 10'b0000000000;
    pxcRom[5579] <= 10'b0000000000;
    pxcRom[5580] <= 10'b0000000000;
    pxcRom[5581] <= 10'b0000000000;
    pxcRom[5582] <= 10'b0000000000;
    pxcRom[5583] <= 10'b0000000000;
    pxcRom[5584] <= 10'b0000000000;
    pxcRom[5585] <= 10'b0000000000;
    pxcRom[5586] <= 10'b0000000000;
    pxcRom[5587] <= 10'b0000000000;
    pxcRom[5588] <= 10'b0000000000;
    pxcRom[5589] <= 10'b0000000000;
    pxcRom[5590] <= 10'b0000000000;
    pxcRom[5591] <= 10'b0000000000;
    pxcRom[5592] <= 10'b0000000000;
    pxcRom[5593] <= 10'b0000000000;
    pxcRom[5594] <= 10'b0000000000;
    pxcRom[5595] <= 10'b0000000000;
    pxcRom[5596] <= 10'b0000000000;
    pxcRom[5597] <= 10'b0000000000;
    pxcRom[5598] <= 10'b0000000000;
    pxcRom[5599] <= 10'b0000000000;
    pxcRom[5600] <= 10'b0000000000;
    pxcRom[5601] <= 10'b0000000000;
    pxcRom[5602] <= 10'b0000000000;
    pxcRom[5603] <= 10'b0000000000;
    pxcRom[5604] <= 10'b0000000000;
    pxcRom[5605] <= 10'b0000000000;
    pxcRom[5606] <= 10'b0000000000;
    pxcRom[5607] <= 10'b0000000000;
    pxcRom[5608] <= 10'b0000000000;
    pxcRom[5609] <= 10'b0000000000;
    pxcRom[5610] <= 10'b0000000000;
    pxcRom[5611] <= 10'b0000000000;
    pxcRom[5612] <= 10'b0000000000;
    pxcRom[5613] <= 10'b0000000000;
    pxcRom[5614] <= 10'b0000000000;
    pxcRom[5615] <= 10'b0000000000;
    pxcRom[5616] <= 10'b0000000000;
    pxcRom[5617] <= 10'b0000000000;
    pxcRom[5618] <= 10'b0000000000;
    pxcRom[5619] <= 10'b0000000000;
    pxcRom[5620] <= 10'b0000000000;
    pxcRom[5621] <= 10'b0000000000;
    pxcRom[5622] <= 10'b0000000000;
    pxcRom[5623] <= 10'b0000000000;
    pxcRom[5624] <= 10'b0000000000;
    pxcRom[5625] <= 10'b0000000000;
    pxcRom[5626] <= 10'b0000000000;
    pxcRom[5627] <= 10'b0000000000;
    pxcRom[5628] <= 10'b0000000000;
    pxcRom[5629] <= 10'b0000000000;
    pxcRom[5630] <= 10'b0000000000;
    pxcRom[5631] <= 10'b0000000000;
    pxcRom[5632] <= 10'b0000000000;
    pxcRom[5633] <= 10'b0000000000;
    pxcRom[5634] <= 10'b0000000000;
    pxcRom[5635] <= 10'b0000000000;
    pxcRom[5636] <= 10'b0000000000;
    pxcRom[5637] <= 10'b0000000000;
    pxcRom[5638] <= 10'b0000000000;
    pxcRom[5639] <= 10'b0000000000;
    pxcRom[5640] <= 10'b0000000000;
    pxcRom[5641] <= 10'b0000000000;
    pxcRom[5642] <= 10'b0000000000;
    pxcRom[5643] <= 10'b0000000000;
    pxcRom[5644] <= 10'b0000000000;
    pxcRom[5645] <= 10'b0000000000;
    pxcRom[5646] <= 10'b0000000000;
    pxcRom[5647] <= 10'b0000000000;
    pxcRom[5648] <= 10'b0000000000;
    pxcRom[5649] <= 10'b0000000000;
    pxcRom[5650] <= 10'b0000000000;
    pxcRom[5651] <= 10'b0000000000;
    pxcRom[5652] <= 10'b0000000000;
    pxcRom[5653] <= 10'b0000000000;
    pxcRom[5654] <= 10'b0000000000;
    pxcRom[5655] <= 10'b0000000000;
    pxcRom[5656] <= 10'b0000000000;
    pxcRom[5657] <= 10'b0000000000;
    pxcRom[5658] <= 10'b0000000000;
    pxcRom[5659] <= 10'b0000000000;
    pxcRom[5660] <= 10'b0000000000;
    pxcRom[5661] <= 10'b0000000001;
    pxcRom[5662] <= 10'b0000000010;
    pxcRom[5663] <= 10'b0000000011;
    pxcRom[5664] <= 10'b0000000101;
    pxcRom[5665] <= 10'b0000000111;
    pxcRom[5666] <= 10'b0000001001;
    pxcRom[5667] <= 10'b0000001010;
    pxcRom[5668] <= 10'b0000001011;
    pxcRom[5669] <= 10'b0000001011;
    pxcRom[5670] <= 10'b0000001011;
    pxcRom[5671] <= 10'b0000001011;
    pxcRom[5672] <= 10'b0000001011;
    pxcRom[5673] <= 10'b0000001010;
    pxcRom[5674] <= 10'b0000001000;
    pxcRom[5675] <= 10'b0000000110;
    pxcRom[5676] <= 10'b0000000011;
    pxcRom[5677] <= 10'b0000000010;
    pxcRom[5678] <= 10'b0000000001;
    pxcRom[5679] <= 10'b0000000000;
    pxcRom[5680] <= 10'b0000000000;
    pxcRom[5681] <= 10'b0000000000;
    pxcRom[5682] <= 10'b0000000000;
    pxcRom[5683] <= 10'b0000000000;
    pxcRom[5684] <= 10'b0000000000;
    pxcRom[5685] <= 10'b0000000000;
    pxcRom[5686] <= 10'b0000000000;
    pxcRom[5687] <= 10'b0000000001;
    pxcRom[5688] <= 10'b0000000011;
    pxcRom[5689] <= 10'b0000000110;
    pxcRom[5690] <= 10'b0000001011;
    pxcRom[5691] <= 10'b0000010001;
    pxcRom[5692] <= 10'b0000011000;
    pxcRom[5693] <= 10'b0000100000;
    pxcRom[5694] <= 10'b0000100111;
    pxcRom[5695] <= 10'b0000101110;
    pxcRom[5696] <= 10'b0000110010;
    pxcRom[5697] <= 10'b0000110110;
    pxcRom[5698] <= 10'b0000111001;
    pxcRom[5699] <= 10'b0000111010;
    pxcRom[5700] <= 10'b0000111010;
    pxcRom[5701] <= 10'b0000110111;
    pxcRom[5702] <= 10'b0000101111;
    pxcRom[5703] <= 10'b0000100011;
    pxcRom[5704] <= 10'b0000010111;
    pxcRom[5705] <= 10'b0000001101;
    pxcRom[5706] <= 10'b0000000110;
    pxcRom[5707] <= 10'b0000000010;
    pxcRom[5708] <= 10'b0000000000;
    pxcRom[5709] <= 10'b0000000000;
    pxcRom[5710] <= 10'b0000000000;
    pxcRom[5711] <= 10'b0000000000;
    pxcRom[5712] <= 10'b0000000000;
    pxcRom[5713] <= 10'b0000000000;
    pxcRom[5714] <= 10'b0000000001;
    pxcRom[5715] <= 10'b0000000011;
    pxcRom[5716] <= 10'b0000000111;
    pxcRom[5717] <= 10'b0000001101;
    pxcRom[5718] <= 10'b0000010110;
    pxcRom[5719] <= 10'b0000100011;
    pxcRom[5720] <= 10'b0000110001;
    pxcRom[5721] <= 10'b0001000010;
    pxcRom[5722] <= 10'b0001010100;
    pxcRom[5723] <= 10'b0001100101;
    pxcRom[5724] <= 10'b0001110001;
    pxcRom[5725] <= 10'b0001110101;
    pxcRom[5726] <= 10'b0001111001;
    pxcRom[5727] <= 10'b0001111011;
    pxcRom[5728] <= 10'b0001111011;
    pxcRom[5729] <= 10'b0001110010;
    pxcRom[5730] <= 10'b0001011101;
    pxcRom[5731] <= 10'b0001000011;
    pxcRom[5732] <= 10'b0000101001;
    pxcRom[5733] <= 10'b0000010110;
    pxcRom[5734] <= 10'b0000001010;
    pxcRom[5735] <= 10'b0000000100;
    pxcRom[5736] <= 10'b0000000001;
    pxcRom[5737] <= 10'b0000000000;
    pxcRom[5738] <= 10'b0000000000;
    pxcRom[5739] <= 10'b0000000000;
    pxcRom[5740] <= 10'b0000000000;
    pxcRom[5741] <= 10'b0000000000;
    pxcRom[5742] <= 10'b0000000001;
    pxcRom[5743] <= 10'b0000000100;
    pxcRom[5744] <= 10'b0000001001;
    pxcRom[5745] <= 10'b0000010010;
    pxcRom[5746] <= 10'b0000011101;
    pxcRom[5747] <= 10'b0000101100;
    pxcRom[5748] <= 10'b0001000000;
    pxcRom[5749] <= 10'b0001010110;
    pxcRom[5750] <= 10'b0001101011;
    pxcRom[5751] <= 10'b0001110111;
    pxcRom[5752] <= 10'b0001111001;
    pxcRom[5753] <= 10'b0001110100;
    pxcRom[5754] <= 10'b0001110010;
    pxcRom[5755] <= 10'b0001111001;
    pxcRom[5756] <= 10'b0010000111;
    pxcRom[5757] <= 10'b0010010000;
    pxcRom[5758] <= 10'b0001111011;
    pxcRom[5759] <= 10'b0001010101;
    pxcRom[5760] <= 10'b0000110010;
    pxcRom[5761] <= 10'b0000011010;
    pxcRom[5762] <= 10'b0000001100;
    pxcRom[5763] <= 10'b0000000100;
    pxcRom[5764] <= 10'b0000000000;
    pxcRom[5765] <= 10'b0000000000;
    pxcRom[5766] <= 10'b0000000000;
    pxcRom[5767] <= 10'b0000000000;
    pxcRom[5768] <= 10'b0000000000;
    pxcRom[5769] <= 10'b0000000000;
    pxcRom[5770] <= 10'b0000000001;
    pxcRom[5771] <= 10'b0000000100;
    pxcRom[5772] <= 10'b0000001001;
    pxcRom[5773] <= 10'b0000010001;
    pxcRom[5774] <= 10'b0000011100;
    pxcRom[5775] <= 10'b0000101001;
    pxcRom[5776] <= 10'b0000111000;
    pxcRom[5777] <= 10'b0001000111;
    pxcRom[5778] <= 10'b0001001100;
    pxcRom[5779] <= 10'b0001001000;
    pxcRom[5780] <= 10'b0001000001;
    pxcRom[5781] <= 10'b0000111010;
    pxcRom[5782] <= 10'b0000111001;
    pxcRom[5783] <= 10'b0000111111;
    pxcRom[5784] <= 10'b0001010001;
    pxcRom[5785] <= 10'b0001101111;
    pxcRom[5786] <= 10'b0001111001;
    pxcRom[5787] <= 10'b0001011000;
    pxcRom[5788] <= 10'b0000110010;
    pxcRom[5789] <= 10'b0000011001;
    pxcRom[5790] <= 10'b0000001010;
    pxcRom[5791] <= 10'b0000000011;
    pxcRom[5792] <= 10'b0000000000;
    pxcRom[5793] <= 10'b0000000000;
    pxcRom[5794] <= 10'b0000000000;
    pxcRom[5795] <= 10'b0000000000;
    pxcRom[5796] <= 10'b0000000000;
    pxcRom[5797] <= 10'b0000000000;
    pxcRom[5798] <= 10'b0000000001;
    pxcRom[5799] <= 10'b0000000011;
    pxcRom[5800] <= 10'b0000000111;
    pxcRom[5801] <= 10'b0000001100;
    pxcRom[5802] <= 10'b0000010101;
    pxcRom[5803] <= 10'b0000011110;
    pxcRom[5804] <= 10'b0000101000;
    pxcRom[5805] <= 10'b0000101101;
    pxcRom[5806] <= 10'b0000101010;
    pxcRom[5807] <= 10'b0000100100;
    pxcRom[5808] <= 10'b0000011100;
    pxcRom[5809] <= 10'b0000010111;
    pxcRom[5810] <= 10'b0000010110;
    pxcRom[5811] <= 10'b0000011110;
    pxcRom[5812] <= 10'b0000110110;
    pxcRom[5813] <= 10'b0001011110;
    pxcRom[5814] <= 10'b0001110001;
    pxcRom[5815] <= 10'b0001010000;
    pxcRom[5816] <= 10'b0000101100;
    pxcRom[5817] <= 10'b0000010100;
    pxcRom[5818] <= 10'b0000001000;
    pxcRom[5819] <= 10'b0000000010;
    pxcRom[5820] <= 10'b0000000000;
    pxcRom[5821] <= 10'b0000000000;
    pxcRom[5822] <= 10'b0000000000;
    pxcRom[5823] <= 10'b0000000000;
    pxcRom[5824] <= 10'b0000000000;
    pxcRom[5825] <= 10'b0000000000;
    pxcRom[5826] <= 10'b0000000000;
    pxcRom[5827] <= 10'b0000000010;
    pxcRom[5828] <= 10'b0000000101;
    pxcRom[5829] <= 10'b0000001000;
    pxcRom[5830] <= 10'b0000001110;
    pxcRom[5831] <= 10'b0000010101;
    pxcRom[5832] <= 10'b0000011010;
    pxcRom[5833] <= 10'b0000011011;
    pxcRom[5834] <= 10'b0000010111;
    pxcRom[5835] <= 10'b0000010000;
    pxcRom[5836] <= 10'b0000001010;
    pxcRom[5837] <= 10'b0000000111;
    pxcRom[5838] <= 10'b0000001010;
    pxcRom[5839] <= 10'b0000010110;
    pxcRom[5840] <= 10'b0000110101;
    pxcRom[5841] <= 10'b0001100100;
    pxcRom[5842] <= 10'b0001101101;
    pxcRom[5843] <= 10'b0001000101;
    pxcRom[5844] <= 10'b0000100011;
    pxcRom[5845] <= 10'b0000001110;
    pxcRom[5846] <= 10'b0000000101;
    pxcRom[5847] <= 10'b0000000001;
    pxcRom[5848] <= 10'b0000000000;
    pxcRom[5849] <= 10'b0000000000;
    pxcRom[5850] <= 10'b0000000000;
    pxcRom[5851] <= 10'b0000000000;
    pxcRom[5852] <= 10'b0000000000;
    pxcRom[5853] <= 10'b0000000000;
    pxcRom[5854] <= 10'b0000000000;
    pxcRom[5855] <= 10'b0000000001;
    pxcRom[5856] <= 10'b0000000011;
    pxcRom[5857] <= 10'b0000000110;
    pxcRom[5858] <= 10'b0000001001;
    pxcRom[5859] <= 10'b0000001110;
    pxcRom[5860] <= 10'b0000010001;
    pxcRom[5861] <= 10'b0000010001;
    pxcRom[5862] <= 10'b0000001101;
    pxcRom[5863] <= 10'b0000000111;
    pxcRom[5864] <= 10'b0000000011;
    pxcRom[5865] <= 10'b0000000011;
    pxcRom[5866] <= 10'b0000001001;
    pxcRom[5867] <= 10'b0000011101;
    pxcRom[5868] <= 10'b0001000110;
    pxcRom[5869] <= 10'b0001110010;
    pxcRom[5870] <= 10'b0001100100;
    pxcRom[5871] <= 10'b0000111001;
    pxcRom[5872] <= 10'b0000011010;
    pxcRom[5873] <= 10'b0000001010;
    pxcRom[5874] <= 10'b0000000011;
    pxcRom[5875] <= 10'b0000000001;
    pxcRom[5876] <= 10'b0000000000;
    pxcRom[5877] <= 10'b0000000000;
    pxcRom[5878] <= 10'b0000000000;
    pxcRom[5879] <= 10'b0000000000;
    pxcRom[5880] <= 10'b0000000000;
    pxcRom[5881] <= 10'b0000000000;
    pxcRom[5882] <= 10'b0000000000;
    pxcRom[5883] <= 10'b0000000000;
    pxcRom[5884] <= 10'b0000000010;
    pxcRom[5885] <= 10'b0000000100;
    pxcRom[5886] <= 10'b0000000110;
    pxcRom[5887] <= 10'b0000001001;
    pxcRom[5888] <= 10'b0000001011;
    pxcRom[5889] <= 10'b0000001010;
    pxcRom[5890] <= 10'b0000000111;
    pxcRom[5891] <= 10'b0000000100;
    pxcRom[5892] <= 10'b0000000011;
    pxcRom[5893] <= 10'b0000000101;
    pxcRom[5894] <= 10'b0000001111;
    pxcRom[5895] <= 10'b0000101101;
    pxcRom[5896] <= 10'b0001011110;
    pxcRom[5897] <= 10'b0001111011;
    pxcRom[5898] <= 10'b0001011010;
    pxcRom[5899] <= 10'b0000101100;
    pxcRom[5900] <= 10'b0000010010;
    pxcRom[5901] <= 10'b0000000111;
    pxcRom[5902] <= 10'b0000000011;
    pxcRom[5903] <= 10'b0000000001;
    pxcRom[5904] <= 10'b0000000000;
    pxcRom[5905] <= 10'b0000000000;
    pxcRom[5906] <= 10'b0000000000;
    pxcRom[5907] <= 10'b0000000000;
    pxcRom[5908] <= 10'b0000000000;
    pxcRom[5909] <= 10'b0000000000;
    pxcRom[5910] <= 10'b0000000000;
    pxcRom[5911] <= 10'b0000000000;
    pxcRom[5912] <= 10'b0000000001;
    pxcRom[5913] <= 10'b0000000010;
    pxcRom[5914] <= 10'b0000000100;
    pxcRom[5915] <= 10'b0000000110;
    pxcRom[5916] <= 10'b0000000111;
    pxcRom[5917] <= 10'b0000000111;
    pxcRom[5918] <= 10'b0000000110;
    pxcRom[5919] <= 10'b0000000101;
    pxcRom[5920] <= 10'b0000000101;
    pxcRom[5921] <= 10'b0000001010;
    pxcRom[5922] <= 10'b0000011101;
    pxcRom[5923] <= 10'b0001000100;
    pxcRom[5924] <= 10'b0001110101;
    pxcRom[5925] <= 10'b0001111000;
    pxcRom[5926] <= 10'b0001000110;
    pxcRom[5927] <= 10'b0000100000;
    pxcRom[5928] <= 10'b0000001110;
    pxcRom[5929] <= 10'b0000000110;
    pxcRom[5930] <= 10'b0000000011;
    pxcRom[5931] <= 10'b0000000001;
    pxcRom[5932] <= 10'b0000000000;
    pxcRom[5933] <= 10'b0000000000;
    pxcRom[5934] <= 10'b0000000000;
    pxcRom[5935] <= 10'b0000000000;
    pxcRom[5936] <= 10'b0000000000;
    pxcRom[5937] <= 10'b0000000000;
    pxcRom[5938] <= 10'b0000000000;
    pxcRom[5939] <= 10'b0000000000;
    pxcRom[5940] <= 10'b0000000000;
    pxcRom[5941] <= 10'b0000000001;
    pxcRom[5942] <= 10'b0000000011;
    pxcRom[5943] <= 10'b0000000100;
    pxcRom[5944] <= 10'b0000000101;
    pxcRom[5945] <= 10'b0000000101;
    pxcRom[5946] <= 10'b0000000110;
    pxcRom[5947] <= 10'b0000000110;
    pxcRom[5948] <= 10'b0000001001;
    pxcRom[5949] <= 10'b0000010100;
    pxcRom[5950] <= 10'b0000110000;
    pxcRom[5951] <= 10'b0001011010;
    pxcRom[5952] <= 10'b0001111110;
    pxcRom[5953] <= 10'b0001100000;
    pxcRom[5954] <= 10'b0000110001;
    pxcRom[5955] <= 10'b0000010110;
    pxcRom[5956] <= 10'b0000001001;
    pxcRom[5957] <= 10'b0000000100;
    pxcRom[5958] <= 10'b0000000010;
    pxcRom[5959] <= 10'b0000000001;
    pxcRom[5960] <= 10'b0000000000;
    pxcRom[5961] <= 10'b0000000000;
    pxcRom[5962] <= 10'b0000000000;
    pxcRom[5963] <= 10'b0000000000;
    pxcRom[5964] <= 10'b0000000000;
    pxcRom[5965] <= 10'b0000000000;
    pxcRom[5966] <= 10'b0000000000;
    pxcRom[5967] <= 10'b0000000000;
    pxcRom[5968] <= 10'b0000000000;
    pxcRom[5969] <= 10'b0000000001;
    pxcRom[5970] <= 10'b0000000001;
    pxcRom[5971] <= 10'b0000000010;
    pxcRom[5972] <= 10'b0000000011;
    pxcRom[5973] <= 10'b0000000100;
    pxcRom[5974] <= 10'b0000000101;
    pxcRom[5975] <= 10'b0000001000;
    pxcRom[5976] <= 10'b0000001110;
    pxcRom[5977] <= 10'b0000100001;
    pxcRom[5978] <= 10'b0001000011;
    pxcRom[5979] <= 10'b0001101011;
    pxcRom[5980] <= 10'b0001101111;
    pxcRom[5981] <= 10'b0001000010;
    pxcRom[5982] <= 10'b0000100001;
    pxcRom[5983] <= 10'b0000001110;
    pxcRom[5984] <= 10'b0000000110;
    pxcRom[5985] <= 10'b0000000011;
    pxcRom[5986] <= 10'b0000000001;
    pxcRom[5987] <= 10'b0000000000;
    pxcRom[5988] <= 10'b0000000000;
    pxcRom[5989] <= 10'b0000000000;
    pxcRom[5990] <= 10'b0000000000;
    pxcRom[5991] <= 10'b0000000000;
    pxcRom[5992] <= 10'b0000000000;
    pxcRom[5993] <= 10'b0000000000;
    pxcRom[5994] <= 10'b0000000000;
    pxcRom[5995] <= 10'b0000000000;
    pxcRom[5996] <= 10'b0000000000;
    pxcRom[5997] <= 10'b0000000000;
    pxcRom[5998] <= 10'b0000000000;
    pxcRom[5999] <= 10'b0000000001;
    pxcRom[6000] <= 10'b0000000010;
    pxcRom[6001] <= 10'b0000000011;
    pxcRom[6002] <= 10'b0000000101;
    pxcRom[6003] <= 10'b0000001001;
    pxcRom[6004] <= 10'b0000010101;
    pxcRom[6005] <= 10'b0000101110;
    pxcRom[6006] <= 10'b0001010011;
    pxcRom[6007] <= 10'b0001101010;
    pxcRom[6008] <= 10'b0001010010;
    pxcRom[6009] <= 10'b0000101100;
    pxcRom[6010] <= 10'b0000010101;
    pxcRom[6011] <= 10'b0000001001;
    pxcRom[6012] <= 10'b0000000100;
    pxcRom[6013] <= 10'b0000000001;
    pxcRom[6014] <= 10'b0000000000;
    pxcRom[6015] <= 10'b0000000000;
    pxcRom[6016] <= 10'b0000000000;
    pxcRom[6017] <= 10'b0000000000;
    pxcRom[6018] <= 10'b0000000000;
    pxcRom[6019] <= 10'b0000000000;
    pxcRom[6020] <= 10'b0000000000;
    pxcRom[6021] <= 10'b0000000000;
    pxcRom[6022] <= 10'b0000000000;
    pxcRom[6023] <= 10'b0000000000;
    pxcRom[6024] <= 10'b0000000000;
    pxcRom[6025] <= 10'b0000000000;
    pxcRom[6026] <= 10'b0000000000;
    pxcRom[6027] <= 10'b0000000000;
    pxcRom[6028] <= 10'b0000000001;
    pxcRom[6029] <= 10'b0000000010;
    pxcRom[6030] <= 10'b0000000101;
    pxcRom[6031] <= 10'b0000001110;
    pxcRom[6032] <= 10'b0000011111;
    pxcRom[6033] <= 10'b0000111010;
    pxcRom[6034] <= 10'b0001011001;
    pxcRom[6035] <= 10'b0001011000;
    pxcRom[6036] <= 10'b0000111001;
    pxcRom[6037] <= 10'b0000011101;
    pxcRom[6038] <= 10'b0000001101;
    pxcRom[6039] <= 10'b0000000101;
    pxcRom[6040] <= 10'b0000000010;
    pxcRom[6041] <= 10'b0000000000;
    pxcRom[6042] <= 10'b0000000000;
    pxcRom[6043] <= 10'b0000000000;
    pxcRom[6044] <= 10'b0000000000;
    pxcRom[6045] <= 10'b0000000000;
    pxcRom[6046] <= 10'b0000000000;
    pxcRom[6047] <= 10'b0000000000;
    pxcRom[6048] <= 10'b0000000000;
    pxcRom[6049] <= 10'b0000000000;
    pxcRom[6050] <= 10'b0000000000;
    pxcRom[6051] <= 10'b0000000000;
    pxcRom[6052] <= 10'b0000000000;
    pxcRom[6053] <= 10'b0000000000;
    pxcRom[6054] <= 10'b0000000000;
    pxcRom[6055] <= 10'b0000000000;
    pxcRom[6056] <= 10'b0000000001;
    pxcRom[6057] <= 10'b0000000011;
    pxcRom[6058] <= 10'b0000001001;
    pxcRom[6059] <= 10'b0000010101;
    pxcRom[6060] <= 10'b0000101001;
    pxcRom[6061] <= 10'b0001000011;
    pxcRom[6062] <= 10'b0001010011;
    pxcRom[6063] <= 10'b0001000011;
    pxcRom[6064] <= 10'b0000100111;
    pxcRom[6065] <= 10'b0000010100;
    pxcRom[6066] <= 10'b0000001001;
    pxcRom[6067] <= 10'b0000000011;
    pxcRom[6068] <= 10'b0000000001;
    pxcRom[6069] <= 10'b0000000000;
    pxcRom[6070] <= 10'b0000000000;
    pxcRom[6071] <= 10'b0000000000;
    pxcRom[6072] <= 10'b0000000000;
    pxcRom[6073] <= 10'b0000000000;
    pxcRom[6074] <= 10'b0000000000;
    pxcRom[6075] <= 10'b0000000000;
    pxcRom[6076] <= 10'b0000000000;
    pxcRom[6077] <= 10'b0000000000;
    pxcRom[6078] <= 10'b0000000000;
    pxcRom[6079] <= 10'b0000000000;
    pxcRom[6080] <= 10'b0000000000;
    pxcRom[6081] <= 10'b0000000000;
    pxcRom[6082] <= 10'b0000000000;
    pxcRom[6083] <= 10'b0000000001;
    pxcRom[6084] <= 10'b0000000011;
    pxcRom[6085] <= 10'b0000000111;
    pxcRom[6086] <= 10'b0000001111;
    pxcRom[6087] <= 10'b0000011110;
    pxcRom[6088] <= 10'b0000110010;
    pxcRom[6089] <= 10'b0001000100;
    pxcRom[6090] <= 10'b0001000100;
    pxcRom[6091] <= 10'b0000110001;
    pxcRom[6092] <= 10'b0000011110;
    pxcRom[6093] <= 10'b0000010000;
    pxcRom[6094] <= 10'b0000000111;
    pxcRom[6095] <= 10'b0000000011;
    pxcRom[6096] <= 10'b0000000001;
    pxcRom[6097] <= 10'b0000000000;
    pxcRom[6098] <= 10'b0000000000;
    pxcRom[6099] <= 10'b0000000000;
    pxcRom[6100] <= 10'b0000000000;
    pxcRom[6101] <= 10'b0000000000;
    pxcRom[6102] <= 10'b0000000000;
    pxcRom[6103] <= 10'b0000000000;
    pxcRom[6104] <= 10'b0000000000;
    pxcRom[6105] <= 10'b0000000000;
    pxcRom[6106] <= 10'b0000000000;
    pxcRom[6107] <= 10'b0000000000;
    pxcRom[6108] <= 10'b0000000000;
    pxcRom[6109] <= 10'b0000000000;
    pxcRom[6110] <= 10'b0000000000;
    pxcRom[6111] <= 10'b0000000010;
    pxcRom[6112] <= 10'b0000000101;
    pxcRom[6113] <= 10'b0000001100;
    pxcRom[6114] <= 10'b0000010110;
    pxcRom[6115] <= 10'b0000100101;
    pxcRom[6116] <= 10'b0000110110;
    pxcRom[6117] <= 10'b0000111110;
    pxcRom[6118] <= 10'b0000110111;
    pxcRom[6119] <= 10'b0000100111;
    pxcRom[6120] <= 10'b0000011000;
    pxcRom[6121] <= 10'b0000001101;
    pxcRom[6122] <= 10'b0000000110;
    pxcRom[6123] <= 10'b0000000010;
    pxcRom[6124] <= 10'b0000000001;
    pxcRom[6125] <= 10'b0000000000;
    pxcRom[6126] <= 10'b0000000000;
    pxcRom[6127] <= 10'b0000000000;
    pxcRom[6128] <= 10'b0000000000;
    pxcRom[6129] <= 10'b0000000000;
    pxcRom[6130] <= 10'b0000000000;
    pxcRom[6131] <= 10'b0000000000;
    pxcRom[6132] <= 10'b0000000000;
    pxcRom[6133] <= 10'b0000000000;
    pxcRom[6134] <= 10'b0000000000;
    pxcRom[6135] <= 10'b0000000000;
    pxcRom[6136] <= 10'b0000000000;
    pxcRom[6137] <= 10'b0000000000;
    pxcRom[6138] <= 10'b0000000010;
    pxcRom[6139] <= 10'b0000000100;
    pxcRom[6140] <= 10'b0000001001;
    pxcRom[6141] <= 10'b0000010001;
    pxcRom[6142] <= 10'b0000011101;
    pxcRom[6143] <= 10'b0000101010;
    pxcRom[6144] <= 10'b0000110100;
    pxcRom[6145] <= 10'b0000110101;
    pxcRom[6146] <= 10'b0000101100;
    pxcRom[6147] <= 10'b0000011111;
    pxcRom[6148] <= 10'b0000010100;
    pxcRom[6149] <= 10'b0000001011;
    pxcRom[6150] <= 10'b0000000101;
    pxcRom[6151] <= 10'b0000000010;
    pxcRom[6152] <= 10'b0000000001;
    pxcRom[6153] <= 10'b0000000000;
    pxcRom[6154] <= 10'b0000000000;
    pxcRom[6155] <= 10'b0000000000;
    pxcRom[6156] <= 10'b0000000000;
    pxcRom[6157] <= 10'b0000000000;
    pxcRom[6158] <= 10'b0000000000;
    pxcRom[6159] <= 10'b0000000000;
    pxcRom[6160] <= 10'b0000000000;
    pxcRom[6161] <= 10'b0000000000;
    pxcRom[6162] <= 10'b0000000000;
    pxcRom[6163] <= 10'b0000000000;
    pxcRom[6164] <= 10'b0000000000;
    pxcRom[6165] <= 10'b0000000001;
    pxcRom[6166] <= 10'b0000000010;
    pxcRom[6167] <= 10'b0000000110;
    pxcRom[6168] <= 10'b0000001100;
    pxcRom[6169] <= 10'b0000010100;
    pxcRom[6170] <= 10'b0000011111;
    pxcRom[6171] <= 10'b0000101001;
    pxcRom[6172] <= 10'b0000101110;
    pxcRom[6173] <= 10'b0000101100;
    pxcRom[6174] <= 10'b0000100011;
    pxcRom[6175] <= 10'b0000011010;
    pxcRom[6176] <= 10'b0000010001;
    pxcRom[6177] <= 10'b0000001001;
    pxcRom[6178] <= 10'b0000000101;
    pxcRom[6179] <= 10'b0000000010;
    pxcRom[6180] <= 10'b0000000001;
    pxcRom[6181] <= 10'b0000000000;
    pxcRom[6182] <= 10'b0000000000;
    pxcRom[6183] <= 10'b0000000000;
    pxcRom[6184] <= 10'b0000000000;
    pxcRom[6185] <= 10'b0000000000;
    pxcRom[6186] <= 10'b0000000000;
    pxcRom[6187] <= 10'b0000000000;
    pxcRom[6188] <= 10'b0000000000;
    pxcRom[6189] <= 10'b0000000000;
    pxcRom[6190] <= 10'b0000000000;
    pxcRom[6191] <= 10'b0000000000;
    pxcRom[6192] <= 10'b0000000000;
    pxcRom[6193] <= 10'b0000000001;
    pxcRom[6194] <= 10'b0000000011;
    pxcRom[6195] <= 10'b0000000110;
    pxcRom[6196] <= 10'b0000001100;
    pxcRom[6197] <= 10'b0000010100;
    pxcRom[6198] <= 10'b0000011101;
    pxcRom[6199] <= 10'b0000100010;
    pxcRom[6200] <= 10'b0000100100;
    pxcRom[6201] <= 10'b0000100001;
    pxcRom[6202] <= 10'b0000011011;
    pxcRom[6203] <= 10'b0000010100;
    pxcRom[6204] <= 10'b0000001101;
    pxcRom[6205] <= 10'b0000001000;
    pxcRom[6206] <= 10'b0000000100;
    pxcRom[6207] <= 10'b0000000010;
    pxcRom[6208] <= 10'b0000000000;
    pxcRom[6209] <= 10'b0000000000;
    pxcRom[6210] <= 10'b0000000000;
    pxcRom[6211] <= 10'b0000000000;
    pxcRom[6212] <= 10'b0000000000;
    pxcRom[6213] <= 10'b0000000000;
    pxcRom[6214] <= 10'b0000000000;
    pxcRom[6215] <= 10'b0000000000;
    pxcRom[6216] <= 10'b0000000000;
    pxcRom[6217] <= 10'b0000000000;
    pxcRom[6218] <= 10'b0000000000;
    pxcRom[6219] <= 10'b0000000000;
    pxcRom[6220] <= 10'b0000000000;
    pxcRom[6221] <= 10'b0000000000;
    pxcRom[6222] <= 10'b0000000001;
    pxcRom[6223] <= 10'b0000000011;
    pxcRom[6224] <= 10'b0000000111;
    pxcRom[6225] <= 10'b0000001010;
    pxcRom[6226] <= 10'b0000001110;
    pxcRom[6227] <= 10'b0000010001;
    pxcRom[6228] <= 10'b0000010010;
    pxcRom[6229] <= 10'b0000010010;
    pxcRom[6230] <= 10'b0000001111;
    pxcRom[6231] <= 10'b0000001011;
    pxcRom[6232] <= 10'b0000001000;
    pxcRom[6233] <= 10'b0000000101;
    pxcRom[6234] <= 10'b0000000010;
    pxcRom[6235] <= 10'b0000000001;
    pxcRom[6236] <= 10'b0000000000;
    pxcRom[6237] <= 10'b0000000000;
    pxcRom[6238] <= 10'b0000000000;
    pxcRom[6239] <= 10'b0000000000;
    pxcRom[6240] <= 10'b0000000000;
    pxcRom[6241] <= 10'b0000000000;
    pxcRom[6242] <= 10'b0000000000;
    pxcRom[6243] <= 10'b0000000000;
    pxcRom[6244] <= 10'b0000000000;
    pxcRom[6245] <= 10'b0000000000;
    pxcRom[6246] <= 10'b0000000000;
    pxcRom[6247] <= 10'b0000000000;
    pxcRom[6248] <= 10'b0000000000;
    pxcRom[6249] <= 10'b0000000000;
    pxcRom[6250] <= 10'b0000000000;
    pxcRom[6251] <= 10'b0000000000;
    pxcRom[6252] <= 10'b0000000000;
    pxcRom[6253] <= 10'b0000000000;
    pxcRom[6254] <= 10'b0000000001;
    pxcRom[6255] <= 10'b0000000001;
    pxcRom[6256] <= 10'b0000000001;
    pxcRom[6257] <= 10'b0000000010;
    pxcRom[6258] <= 10'b0000000010;
    pxcRom[6259] <= 10'b0000000010;
    pxcRom[6260] <= 10'b0000000001;
    pxcRom[6261] <= 10'b0000000001;
    pxcRom[6262] <= 10'b0000000000;
    pxcRom[6263] <= 10'b0000000000;
    pxcRom[6264] <= 10'b0000000000;
    pxcRom[6265] <= 10'b0000000000;
    pxcRom[6266] <= 10'b0000000000;
    pxcRom[6267] <= 10'b0000000000;
    pxcRom[6268] <= 10'b0000000000;
    pxcRom[6269] <= 10'b0000000000;
    pxcRom[6270] <= 10'b0000000000;
    pxcRom[6271] <= 10'b0000000000;
    pxcRom[6272] <= 10'b0000000000;
    pxcRom[6273] <= 10'b0000000000;
    pxcRom[6274] <= 10'b0000000000;
    pxcRom[6275] <= 10'b0000000000;
    pxcRom[6276] <= 10'b0000000000;
    pxcRom[6277] <= 10'b0000000000;
    pxcRom[6278] <= 10'b0000000000;
    pxcRom[6279] <= 10'b0000000000;
    pxcRom[6280] <= 10'b0000000000;
    pxcRom[6281] <= 10'b0000000000;
    pxcRom[6282] <= 10'b0000000000;
    pxcRom[6283] <= 10'b0000000000;
    pxcRom[6284] <= 10'b0000000000;
    pxcRom[6285] <= 10'b0000000000;
    pxcRom[6286] <= 10'b0000000000;
    pxcRom[6287] <= 10'b0000000000;
    pxcRom[6288] <= 10'b0000000000;
    pxcRom[6289] <= 10'b0000000000;
    pxcRom[6290] <= 10'b0000000000;
    pxcRom[6291] <= 10'b0000000000;
    pxcRom[6292] <= 10'b0000000000;
    pxcRom[6293] <= 10'b0000000000;
    pxcRom[6294] <= 10'b0000000000;
    pxcRom[6295] <= 10'b0000000000;
    pxcRom[6296] <= 10'b0000000000;
    pxcRom[6297] <= 10'b0000000000;
    pxcRom[6298] <= 10'b0000000000;
    pxcRom[6299] <= 10'b0000000000;
    pxcRom[6300] <= 10'b0000000000;
    pxcRom[6301] <= 10'b0000000000;
    pxcRom[6302] <= 10'b0000000000;
    pxcRom[6303] <= 10'b0000000000;
    pxcRom[6304] <= 10'b0000000000;
    pxcRom[6305] <= 10'b0000000000;
    pxcRom[6306] <= 10'b0000000000;
    pxcRom[6307] <= 10'b0000000000;
    pxcRom[6308] <= 10'b0000000000;
    pxcRom[6309] <= 10'b0000000000;
    pxcRom[6310] <= 10'b0000000000;
    pxcRom[6311] <= 10'b0000000000;
    pxcRom[6312] <= 10'b0000000000;
    pxcRom[6313] <= 10'b0000000000;
    pxcRom[6314] <= 10'b0000000000;
    pxcRom[6315] <= 10'b0000000000;
    pxcRom[6316] <= 10'b0000000000;
    pxcRom[6317] <= 10'b0000000000;
    pxcRom[6318] <= 10'b0000000000;
    pxcRom[6319] <= 10'b0000000000;
    pxcRom[6320] <= 10'b0000000000;
    pxcRom[6321] <= 10'b0000000000;
    pxcRom[6322] <= 10'b0000000000;
    pxcRom[6323] <= 10'b0000000000;
    pxcRom[6324] <= 10'b0000000000;
    pxcRom[6325] <= 10'b0000000000;
    pxcRom[6326] <= 10'b0000000000;
    pxcRom[6327] <= 10'b0000000000;
    pxcRom[6328] <= 10'b0000000000;
    pxcRom[6329] <= 10'b0000000000;
    pxcRom[6330] <= 10'b0000000000;
    pxcRom[6331] <= 10'b0000000000;
    pxcRom[6332] <= 10'b0000000000;
    pxcRom[6333] <= 10'b0000000000;
    pxcRom[6334] <= 10'b0000000000;
    pxcRom[6335] <= 10'b0000000000;
    pxcRom[6336] <= 10'b0000000000;
    pxcRom[6337] <= 10'b0000000000;
    pxcRom[6338] <= 10'b0000000000;
    pxcRom[6339] <= 10'b0000000000;
    pxcRom[6340] <= 10'b0000000000;
    pxcRom[6341] <= 10'b0000000000;
    pxcRom[6342] <= 10'b0000000000;
    pxcRom[6343] <= 10'b0000000000;
    pxcRom[6344] <= 10'b0000000000;
    pxcRom[6345] <= 10'b0000000000;
    pxcRom[6346] <= 10'b0000000000;
    pxcRom[6347] <= 10'b0000000000;
    pxcRom[6348] <= 10'b0000000000;
    pxcRom[6349] <= 10'b0000000000;
    pxcRom[6350] <= 10'b0000000000;
    pxcRom[6351] <= 10'b0000000000;
    pxcRom[6352] <= 10'b0000000000;
    pxcRom[6353] <= 10'b0000000000;
    pxcRom[6354] <= 10'b0000000000;
    pxcRom[6355] <= 10'b0000000000;
    pxcRom[6356] <= 10'b0000000000;
    pxcRom[6357] <= 10'b0000000000;
    pxcRom[6358] <= 10'b0000000000;
    pxcRom[6359] <= 10'b0000000000;
    pxcRom[6360] <= 10'b0000000000;
    pxcRom[6361] <= 10'b0000000000;
    pxcRom[6362] <= 10'b0000000000;
    pxcRom[6363] <= 10'b0000000000;
    pxcRom[6364] <= 10'b0000000000;
    pxcRom[6365] <= 10'b0000000000;
    pxcRom[6366] <= 10'b0000000000;
    pxcRom[6367] <= 10'b0000000000;
    pxcRom[6368] <= 10'b0000000000;
    pxcRom[6369] <= 10'b0000000000;
    pxcRom[6370] <= 10'b0000000000;
    pxcRom[6371] <= 10'b0000000000;
    pxcRom[6372] <= 10'b0000000000;
    pxcRom[6373] <= 10'b0000000000;
    pxcRom[6374] <= 10'b0000000000;
    pxcRom[6375] <= 10'b0000000000;
    pxcRom[6376] <= 10'b0000000000;
    pxcRom[6377] <= 10'b0000000000;
    pxcRom[6378] <= 10'b0000000000;
    pxcRom[6379] <= 10'b0000000000;
    pxcRom[6380] <= 10'b0000000000;
    pxcRom[6381] <= 10'b0000000000;
    pxcRom[6382] <= 10'b0000000000;
    pxcRom[6383] <= 10'b0000000000;
    pxcRom[6384] <= 10'b0000000000;
    pxcRom[6385] <= 10'b0000000000;
    pxcRom[6386] <= 10'b0000000000;
    pxcRom[6387] <= 10'b0000000000;
    pxcRom[6388] <= 10'b0000000000;
    pxcRom[6389] <= 10'b0000000000;
    pxcRom[6390] <= 10'b0000000000;
    pxcRom[6391] <= 10'b0000000000;
    pxcRom[6392] <= 10'b0000000000;
    pxcRom[6393] <= 10'b0000000000;
    pxcRom[6394] <= 10'b0000000001;
    pxcRom[6395] <= 10'b0000000011;
    pxcRom[6396] <= 10'b0000000101;
    pxcRom[6397] <= 10'b0000001000;
    pxcRom[6398] <= 10'b0000001011;
    pxcRom[6399] <= 10'b0000001101;
    pxcRom[6400] <= 10'b0000001101;
    pxcRom[6401] <= 10'b0000001100;
    pxcRom[6402] <= 10'b0000001001;
    pxcRom[6403] <= 10'b0000000110;
    pxcRom[6404] <= 10'b0000000100;
    pxcRom[6405] <= 10'b0000000010;
    pxcRom[6406] <= 10'b0000000001;
    pxcRom[6407] <= 10'b0000000000;
    pxcRom[6408] <= 10'b0000000000;
    pxcRom[6409] <= 10'b0000000000;
    pxcRom[6410] <= 10'b0000000000;
    pxcRom[6411] <= 10'b0000000000;
    pxcRom[6412] <= 10'b0000000000;
    pxcRom[6413] <= 10'b0000000000;
    pxcRom[6414] <= 10'b0000000000;
    pxcRom[6415] <= 10'b0000000000;
    pxcRom[6416] <= 10'b0000000000;
    pxcRom[6417] <= 10'b0000000000;
    pxcRom[6418] <= 10'b0000000000;
    pxcRom[6419] <= 10'b0000000000;
    pxcRom[6420] <= 10'b0000000010;
    pxcRom[6421] <= 10'b0000000101;
    pxcRom[6422] <= 10'b0000001010;
    pxcRom[6423] <= 10'b0000010010;
    pxcRom[6424] <= 10'b0000011111;
    pxcRom[6425] <= 10'b0000101101;
    pxcRom[6426] <= 10'b0000111110;
    pxcRom[6427] <= 10'b0001001010;
    pxcRom[6428] <= 10'b0001001101;
    pxcRom[6429] <= 10'b0001000100;
    pxcRom[6430] <= 10'b0000110011;
    pxcRom[6431] <= 10'b0000100011;
    pxcRom[6432] <= 10'b0000010111;
    pxcRom[6433] <= 10'b0000001101;
    pxcRom[6434] <= 10'b0000000111;
    pxcRom[6435] <= 10'b0000000011;
    pxcRom[6436] <= 10'b0000000001;
    pxcRom[6437] <= 10'b0000000000;
    pxcRom[6438] <= 10'b0000000000;
    pxcRom[6439] <= 10'b0000000000;
    pxcRom[6440] <= 10'b0000000000;
    pxcRom[6441] <= 10'b0000000000;
    pxcRom[6442] <= 10'b0000000000;
    pxcRom[6443] <= 10'b0000000000;
    pxcRom[6444] <= 10'b0000000000;
    pxcRom[6445] <= 10'b0000000000;
    pxcRom[6446] <= 10'b0000000001;
    pxcRom[6447] <= 10'b0000000011;
    pxcRom[6448] <= 10'b0000000111;
    pxcRom[6449] <= 10'b0000001110;
    pxcRom[6450] <= 10'b0000011010;
    pxcRom[6451] <= 10'b0000101100;
    pxcRom[6452] <= 10'b0001000011;
    pxcRom[6453] <= 10'b0001011101;
    pxcRom[6454] <= 10'b0001110011;
    pxcRom[6455] <= 10'b0001111111;
    pxcRom[6456] <= 10'b0001111101;
    pxcRom[6457] <= 10'b0001101100;
    pxcRom[6458] <= 10'b0001010110;
    pxcRom[6459] <= 10'b0000111101;
    pxcRom[6460] <= 10'b0000101001;
    pxcRom[6461] <= 10'b0000011001;
    pxcRom[6462] <= 10'b0000001110;
    pxcRom[6463] <= 10'b0000001000;
    pxcRom[6464] <= 10'b0000000011;
    pxcRom[6465] <= 10'b0000000001;
    pxcRom[6466] <= 10'b0000000000;
    pxcRom[6467] <= 10'b0000000000;
    pxcRom[6468] <= 10'b0000000000;
    pxcRom[6469] <= 10'b0000000000;
    pxcRom[6470] <= 10'b0000000000;
    pxcRom[6471] <= 10'b0000000000;
    pxcRom[6472] <= 10'b0000000000;
    pxcRom[6473] <= 10'b0000000000;
    pxcRom[6474] <= 10'b0000000010;
    pxcRom[6475] <= 10'b0000000111;
    pxcRom[6476] <= 10'b0000001101;
    pxcRom[6477] <= 10'b0000011001;
    pxcRom[6478] <= 10'b0000101100;
    pxcRom[6479] <= 10'b0001000100;
    pxcRom[6480] <= 10'b0001011100;
    pxcRom[6481] <= 10'b0001101010;
    pxcRom[6482] <= 10'b0001100101;
    pxcRom[6483] <= 10'b0001100000;
    pxcRom[6484] <= 10'b0001011100;
    pxcRom[6485] <= 10'b0001011011;
    pxcRom[6486] <= 10'b0001010110;
    pxcRom[6487] <= 10'b0001001000;
    pxcRom[6488] <= 10'b0000110101;
    pxcRom[6489] <= 10'b0000100010;
    pxcRom[6490] <= 10'b0000010101;
    pxcRom[6491] <= 10'b0000001100;
    pxcRom[6492] <= 10'b0000000101;
    pxcRom[6493] <= 10'b0000000001;
    pxcRom[6494] <= 10'b0000000000;
    pxcRom[6495] <= 10'b0000000000;
    pxcRom[6496] <= 10'b0000000000;
    pxcRom[6497] <= 10'b0000000000;
    pxcRom[6498] <= 10'b0000000000;
    pxcRom[6499] <= 10'b0000000000;
    pxcRom[6500] <= 10'b0000000000;
    pxcRom[6501] <= 10'b0000000001;
    pxcRom[6502] <= 10'b0000000100;
    pxcRom[6503] <= 10'b0000001010;
    pxcRom[6504] <= 10'b0000010100;
    pxcRom[6505] <= 10'b0000100101;
    pxcRom[6506] <= 10'b0000111011;
    pxcRom[6507] <= 10'b0001001111;
    pxcRom[6508] <= 10'b0001010101;
    pxcRom[6509] <= 10'b0001001011;
    pxcRom[6510] <= 10'b0000111011;
    pxcRom[6511] <= 10'b0000110001;
    pxcRom[6512] <= 10'b0000110010;
    pxcRom[6513] <= 10'b0000111000;
    pxcRom[6514] <= 10'b0001000011;
    pxcRom[6515] <= 10'b0001000111;
    pxcRom[6516] <= 10'b0000111001;
    pxcRom[6517] <= 10'b0000100111;
    pxcRom[6518] <= 10'b0000011001;
    pxcRom[6519] <= 10'b0000001110;
    pxcRom[6520] <= 10'b0000000111;
    pxcRom[6521] <= 10'b0000000010;
    pxcRom[6522] <= 10'b0000000000;
    pxcRom[6523] <= 10'b0000000000;
    pxcRom[6524] <= 10'b0000000000;
    pxcRom[6525] <= 10'b0000000000;
    pxcRom[6526] <= 10'b0000000000;
    pxcRom[6527] <= 10'b0000000000;
    pxcRom[6528] <= 10'b0000000000;
    pxcRom[6529] <= 10'b0000000010;
    pxcRom[6530] <= 10'b0000000110;
    pxcRom[6531] <= 10'b0000001101;
    pxcRom[6532] <= 10'b0000011001;
    pxcRom[6533] <= 10'b0000101100;
    pxcRom[6534] <= 10'b0001000000;
    pxcRom[6535] <= 10'b0001001011;
    pxcRom[6536] <= 10'b0001000011;
    pxcRom[6537] <= 10'b0000101111;
    pxcRom[6538] <= 10'b0000100001;
    pxcRom[6539] <= 10'b0000011011;
    pxcRom[6540] <= 10'b0000100000;
    pxcRom[6541] <= 10'b0000101110;
    pxcRom[6542] <= 10'b0001000000;
    pxcRom[6543] <= 10'b0001001000;
    pxcRom[6544] <= 10'b0000111011;
    pxcRom[6545] <= 10'b0000101000;
    pxcRom[6546] <= 10'b0000011000;
    pxcRom[6547] <= 10'b0000001101;
    pxcRom[6548] <= 10'b0000000110;
    pxcRom[6549] <= 10'b0000000010;
    pxcRom[6550] <= 10'b0000000000;
    pxcRom[6551] <= 10'b0000000000;
    pxcRom[6552] <= 10'b0000000000;
    pxcRom[6553] <= 10'b0000000000;
    pxcRom[6554] <= 10'b0000000000;
    pxcRom[6555] <= 10'b0000000000;
    pxcRom[6556] <= 10'b0000000000;
    pxcRom[6557] <= 10'b0000000010;
    pxcRom[6558] <= 10'b0000000110;
    pxcRom[6559] <= 10'b0000001110;
    pxcRom[6560] <= 10'b0000011010;
    pxcRom[6561] <= 10'b0000101101;
    pxcRom[6562] <= 10'b0001000001;
    pxcRom[6563] <= 10'b0001000111;
    pxcRom[6564] <= 10'b0000111010;
    pxcRom[6565] <= 10'b0000100110;
    pxcRom[6566] <= 10'b0000011001;
    pxcRom[6567] <= 10'b0000011001;
    pxcRom[6568] <= 10'b0000100011;
    pxcRom[6569] <= 10'b0000110111;
    pxcRom[6570] <= 10'b0001001100;
    pxcRom[6571] <= 10'b0001001001;
    pxcRom[6572] <= 10'b0000110111;
    pxcRom[6573] <= 10'b0000100010;
    pxcRom[6574] <= 10'b0000010100;
    pxcRom[6575] <= 10'b0000001010;
    pxcRom[6576] <= 10'b0000000101;
    pxcRom[6577] <= 10'b0000000001;
    pxcRom[6578] <= 10'b0000000000;
    pxcRom[6579] <= 10'b0000000000;
    pxcRom[6580] <= 10'b0000000000;
    pxcRom[6581] <= 10'b0000000000;
    pxcRom[6582] <= 10'b0000000000;
    pxcRom[6583] <= 10'b0000000000;
    pxcRom[6584] <= 10'b0000000000;
    pxcRom[6585] <= 10'b0000000010;
    pxcRom[6586] <= 10'b0000000110;
    pxcRom[6587] <= 10'b0000001101;
    pxcRom[6588] <= 10'b0000011000;
    pxcRom[6589] <= 10'b0000101011;
    pxcRom[6590] <= 10'b0000111110;
    pxcRom[6591] <= 10'b0001001000;
    pxcRom[6592] <= 10'b0001000000;
    pxcRom[6593] <= 10'b0000101101;
    pxcRom[6594] <= 10'b0000100010;
    pxcRom[6595] <= 10'b0000100111;
    pxcRom[6596] <= 10'b0000111010;
    pxcRom[6597] <= 10'b0001010000;
    pxcRom[6598] <= 10'b0001010101;
    pxcRom[6599] <= 10'b0001000010;
    pxcRom[6600] <= 10'b0000101001;
    pxcRom[6601] <= 10'b0000011000;
    pxcRom[6602] <= 10'b0000001101;
    pxcRom[6603] <= 10'b0000000110;
    pxcRom[6604] <= 10'b0000000011;
    pxcRom[6605] <= 10'b0000000001;
    pxcRom[6606] <= 10'b0000000000;
    pxcRom[6607] <= 10'b0000000000;
    pxcRom[6608] <= 10'b0000000000;
    pxcRom[6609] <= 10'b0000000000;
    pxcRom[6610] <= 10'b0000000000;
    pxcRom[6611] <= 10'b0000000000;
    pxcRom[6612] <= 10'b0000000000;
    pxcRom[6613] <= 10'b0000000001;
    pxcRom[6614] <= 10'b0000000100;
    pxcRom[6615] <= 10'b0000001010;
    pxcRom[6616] <= 10'b0000010100;
    pxcRom[6617] <= 10'b0000100011;
    pxcRom[6618] <= 10'b0000111000;
    pxcRom[6619] <= 10'b0001001100;
    pxcRom[6620] <= 10'b0001010000;
    pxcRom[6621] <= 10'b0001000101;
    pxcRom[6622] <= 10'b0000111101;
    pxcRom[6623] <= 10'b0001001010;
    pxcRom[6624] <= 10'b0001100000;
    pxcRom[6625] <= 10'b0001100011;
    pxcRom[6626] <= 10'b0001001010;
    pxcRom[6627] <= 10'b0000101111;
    pxcRom[6628] <= 10'b0000011011;
    pxcRom[6629] <= 10'b0000001110;
    pxcRom[6630] <= 10'b0000000111;
    pxcRom[6631] <= 10'b0000000011;
    pxcRom[6632] <= 10'b0000000001;
    pxcRom[6633] <= 10'b0000000000;
    pxcRom[6634] <= 10'b0000000000;
    pxcRom[6635] <= 10'b0000000000;
    pxcRom[6636] <= 10'b0000000000;
    pxcRom[6637] <= 10'b0000000000;
    pxcRom[6638] <= 10'b0000000000;
    pxcRom[6639] <= 10'b0000000000;
    pxcRom[6640] <= 10'b0000000000;
    pxcRom[6641] <= 10'b0000000001;
    pxcRom[6642] <= 10'b0000000011;
    pxcRom[6643] <= 10'b0000000111;
    pxcRom[6644] <= 10'b0000001110;
    pxcRom[6645] <= 10'b0000011011;
    pxcRom[6646] <= 10'b0000101101;
    pxcRom[6647] <= 10'b0001001011;
    pxcRom[6648] <= 10'b0001101001;
    pxcRom[6649] <= 10'b0001101111;
    pxcRom[6650] <= 10'b0001101100;
    pxcRom[6651] <= 10'b0001111111;
    pxcRom[6652] <= 10'b0001111110;
    pxcRom[6653] <= 10'b0001011000;
    pxcRom[6654] <= 10'b0000110100;
    pxcRom[6655] <= 10'b0000011100;
    pxcRom[6656] <= 10'b0000001110;
    pxcRom[6657] <= 10'b0000000111;
    pxcRom[6658] <= 10'b0000000011;
    pxcRom[6659] <= 10'b0000000001;
    pxcRom[6660] <= 10'b0000000000;
    pxcRom[6661] <= 10'b0000000000;
    pxcRom[6662] <= 10'b0000000000;
    pxcRom[6663] <= 10'b0000000000;
    pxcRom[6664] <= 10'b0000000000;
    pxcRom[6665] <= 10'b0000000000;
    pxcRom[6666] <= 10'b0000000000;
    pxcRom[6667] <= 10'b0000000000;
    pxcRom[6668] <= 10'b0000000000;
    pxcRom[6669] <= 10'b0000000000;
    pxcRom[6670] <= 10'b0000000001;
    pxcRom[6671] <= 10'b0000000100;
    pxcRom[6672] <= 10'b0000001001;
    pxcRom[6673] <= 10'b0000010011;
    pxcRom[6674] <= 10'b0000100111;
    pxcRom[6675] <= 10'b0001001000;
    pxcRom[6676] <= 10'b0001111011;
    pxcRom[6677] <= 10'b0010011101;
    pxcRom[6678] <= 10'b0010101010;
    pxcRom[6679] <= 10'b0010100100;
    pxcRom[6680] <= 10'b0001110011;
    pxcRom[6681] <= 10'b0001000000;
    pxcRom[6682] <= 10'b0000100000;
    pxcRom[6683] <= 10'b0000010000;
    pxcRom[6684] <= 10'b0000001000;
    pxcRom[6685] <= 10'b0000000100;
    pxcRom[6686] <= 10'b0000000010;
    pxcRom[6687] <= 10'b0000000001;
    pxcRom[6688] <= 10'b0000000000;
    pxcRom[6689] <= 10'b0000000000;
    pxcRom[6690] <= 10'b0000000000;
    pxcRom[6691] <= 10'b0000000000;
    pxcRom[6692] <= 10'b0000000000;
    pxcRom[6693] <= 10'b0000000000;
    pxcRom[6694] <= 10'b0000000000;
    pxcRom[6695] <= 10'b0000000000;
    pxcRom[6696] <= 10'b0000000000;
    pxcRom[6697] <= 10'b0000000000;
    pxcRom[6698] <= 10'b0000000001;
    pxcRom[6699] <= 10'b0000000011;
    pxcRom[6700] <= 10'b0000001000;
    pxcRom[6701] <= 10'b0000010010;
    pxcRom[6702] <= 10'b0000100110;
    pxcRom[6703] <= 10'b0001001100;
    pxcRom[6704] <= 10'b0010000111;
    pxcRom[6705] <= 10'b0010100111;
    pxcRom[6706] <= 10'b0010100100;
    pxcRom[6707] <= 10'b0010000110;
    pxcRom[6708] <= 10'b0001010111;
    pxcRom[6709] <= 10'b0000101110;
    pxcRom[6710] <= 10'b0000011000;
    pxcRom[6711] <= 10'b0000001100;
    pxcRom[6712] <= 10'b0000000111;
    pxcRom[6713] <= 10'b0000000011;
    pxcRom[6714] <= 10'b0000000010;
    pxcRom[6715] <= 10'b0000000001;
    pxcRom[6716] <= 10'b0000000000;
    pxcRom[6717] <= 10'b0000000000;
    pxcRom[6718] <= 10'b0000000000;
    pxcRom[6719] <= 10'b0000000000;
    pxcRom[6720] <= 10'b0000000000;
    pxcRom[6721] <= 10'b0000000000;
    pxcRom[6722] <= 10'b0000000000;
    pxcRom[6723] <= 10'b0000000000;
    pxcRom[6724] <= 10'b0000000000;
    pxcRom[6725] <= 10'b0000000000;
    pxcRom[6726] <= 10'b0000000001;
    pxcRom[6727] <= 10'b0000000100;
    pxcRom[6728] <= 10'b0000001011;
    pxcRom[6729] <= 10'b0000011000;
    pxcRom[6730] <= 10'b0000110001;
    pxcRom[6731] <= 10'b0001011010;
    pxcRom[6732] <= 10'b0010000000;
    pxcRom[6733] <= 10'b0001111110;
    pxcRom[6734] <= 10'b0001101110;
    pxcRom[6735] <= 10'b0001011101;
    pxcRom[6736] <= 10'b0001000010;
    pxcRom[6737] <= 10'b0000101001;
    pxcRom[6738] <= 10'b0000010111;
    pxcRom[6739] <= 10'b0000001101;
    pxcRom[6740] <= 10'b0000000111;
    pxcRom[6741] <= 10'b0000000100;
    pxcRom[6742] <= 10'b0000000010;
    pxcRom[6743] <= 10'b0000000001;
    pxcRom[6744] <= 10'b0000000000;
    pxcRom[6745] <= 10'b0000000000;
    pxcRom[6746] <= 10'b0000000000;
    pxcRom[6747] <= 10'b0000000000;
    pxcRom[6748] <= 10'b0000000000;
    pxcRom[6749] <= 10'b0000000000;
    pxcRom[6750] <= 10'b0000000000;
    pxcRom[6751] <= 10'b0000000000;
    pxcRom[6752] <= 10'b0000000000;
    pxcRom[6753] <= 10'b0000000000;
    pxcRom[6754] <= 10'b0000000011;
    pxcRom[6755] <= 10'b0000001000;
    pxcRom[6756] <= 10'b0000010010;
    pxcRom[6757] <= 10'b0000100101;
    pxcRom[6758] <= 10'b0001000011;
    pxcRom[6759] <= 10'b0001100011;
    pxcRom[6760] <= 10'b0001100101;
    pxcRom[6761] <= 10'b0001010001;
    pxcRom[6762] <= 10'b0001000101;
    pxcRom[6763] <= 10'b0001000001;
    pxcRom[6764] <= 10'b0000111001;
    pxcRom[6765] <= 10'b0000101001;
    pxcRom[6766] <= 10'b0000011011;
    pxcRom[6767] <= 10'b0000010000;
    pxcRom[6768] <= 10'b0000001001;
    pxcRom[6769] <= 10'b0000000101;
    pxcRom[6770] <= 10'b0000000011;
    pxcRom[6771] <= 10'b0000000001;
    pxcRom[6772] <= 10'b0000000000;
    pxcRom[6773] <= 10'b0000000000;
    pxcRom[6774] <= 10'b0000000000;
    pxcRom[6775] <= 10'b0000000000;
    pxcRom[6776] <= 10'b0000000000;
    pxcRom[6777] <= 10'b0000000000;
    pxcRom[6778] <= 10'b0000000000;
    pxcRom[6779] <= 10'b0000000000;
    pxcRom[6780] <= 10'b0000000000;
    pxcRom[6781] <= 10'b0000000001;
    pxcRom[6782] <= 10'b0000000101;
    pxcRom[6783] <= 10'b0000001101;
    pxcRom[6784] <= 10'b0000011101;
    pxcRom[6785] <= 10'b0000110011;
    pxcRom[6786] <= 10'b0001001111;
    pxcRom[6787] <= 10'b0001010111;
    pxcRom[6788] <= 10'b0001000101;
    pxcRom[6789] <= 10'b0000110011;
    pxcRom[6790] <= 10'b0000101110;
    pxcRom[6791] <= 10'b0000110101;
    pxcRom[6792] <= 10'b0000110101;
    pxcRom[6793] <= 10'b0000101010;
    pxcRom[6794] <= 10'b0000011110;
    pxcRom[6795] <= 10'b0000010011;
    pxcRom[6796] <= 10'b0000001011;
    pxcRom[6797] <= 10'b0000000110;
    pxcRom[6798] <= 10'b0000000011;
    pxcRom[6799] <= 10'b0000000010;
    pxcRom[6800] <= 10'b0000000000;
    pxcRom[6801] <= 10'b0000000000;
    pxcRom[6802] <= 10'b0000000000;
    pxcRom[6803] <= 10'b0000000000;
    pxcRom[6804] <= 10'b0000000000;
    pxcRom[6805] <= 10'b0000000000;
    pxcRom[6806] <= 10'b0000000000;
    pxcRom[6807] <= 10'b0000000000;
    pxcRom[6808] <= 10'b0000000000;
    pxcRom[6809] <= 10'b0000000010;
    pxcRom[6810] <= 10'b0000001000;
    pxcRom[6811] <= 10'b0000010011;
    pxcRom[6812] <= 10'b0000100110;
    pxcRom[6813] <= 10'b0000111101;
    pxcRom[6814] <= 10'b0001001110;
    pxcRom[6815] <= 10'b0001000011;
    pxcRom[6816] <= 10'b0000101111;
    pxcRom[6817] <= 10'b0000100011;
    pxcRom[6818] <= 10'b0000100101;
    pxcRom[6819] <= 10'b0000101111;
    pxcRom[6820] <= 10'b0000110100;
    pxcRom[6821] <= 10'b0000101100;
    pxcRom[6822] <= 10'b0000100001;
    pxcRom[6823] <= 10'b0000010101;
    pxcRom[6824] <= 10'b0000001100;
    pxcRom[6825] <= 10'b0000000111;
    pxcRom[6826] <= 10'b0000000011;
    pxcRom[6827] <= 10'b0000000001;
    pxcRom[6828] <= 10'b0000000000;
    pxcRom[6829] <= 10'b0000000000;
    pxcRom[6830] <= 10'b0000000000;
    pxcRom[6831] <= 10'b0000000000;
    pxcRom[6832] <= 10'b0000000000;
    pxcRom[6833] <= 10'b0000000000;
    pxcRom[6834] <= 10'b0000000000;
    pxcRom[6835] <= 10'b0000000000;
    pxcRom[6836] <= 10'b0000000000;
    pxcRom[6837] <= 10'b0000000011;
    pxcRom[6838] <= 10'b0000001011;
    pxcRom[6839] <= 10'b0000011000;
    pxcRom[6840] <= 10'b0000101010;
    pxcRom[6841] <= 10'b0000111111;
    pxcRom[6842] <= 10'b0001001000;
    pxcRom[6843] <= 10'b0000111010;
    pxcRom[6844] <= 10'b0000101011;
    pxcRom[6845] <= 10'b0000100101;
    pxcRom[6846] <= 10'b0000101011;
    pxcRom[6847] <= 10'b0000110100;
    pxcRom[6848] <= 10'b0000110111;
    pxcRom[6849] <= 10'b0000101111;
    pxcRom[6850] <= 10'b0000100010;
    pxcRom[6851] <= 10'b0000010101;
    pxcRom[6852] <= 10'b0000001100;
    pxcRom[6853] <= 10'b0000000110;
    pxcRom[6854] <= 10'b0000000011;
    pxcRom[6855] <= 10'b0000000001;
    pxcRom[6856] <= 10'b0000000000;
    pxcRom[6857] <= 10'b0000000000;
    pxcRom[6858] <= 10'b0000000000;
    pxcRom[6859] <= 10'b0000000000;
    pxcRom[6860] <= 10'b0000000000;
    pxcRom[6861] <= 10'b0000000000;
    pxcRom[6862] <= 10'b0000000000;
    pxcRom[6863] <= 10'b0000000000;
    pxcRom[6864] <= 10'b0000000000;
    pxcRom[6865] <= 10'b0000000011;
    pxcRom[6866] <= 10'b0000001011;
    pxcRom[6867] <= 10'b0000011001;
    pxcRom[6868] <= 10'b0000101011;
    pxcRom[6869] <= 10'b0000111111;
    pxcRom[6870] <= 10'b0001001100;
    pxcRom[6871] <= 10'b0001001000;
    pxcRom[6872] <= 10'b0001000001;
    pxcRom[6873] <= 10'b0001000000;
    pxcRom[6874] <= 10'b0001000011;
    pxcRom[6875] <= 10'b0001000110;
    pxcRom[6876] <= 10'b0001000000;
    pxcRom[6877] <= 10'b0000110001;
    pxcRom[6878] <= 10'b0000100001;
    pxcRom[6879] <= 10'b0000010100;
    pxcRom[6880] <= 10'b0000001011;
    pxcRom[6881] <= 10'b0000000101;
    pxcRom[6882] <= 10'b0000000010;
    pxcRom[6883] <= 10'b0000000001;
    pxcRom[6884] <= 10'b0000000000;
    pxcRom[6885] <= 10'b0000000000;
    pxcRom[6886] <= 10'b0000000000;
    pxcRom[6887] <= 10'b0000000000;
    pxcRom[6888] <= 10'b0000000000;
    pxcRom[6889] <= 10'b0000000000;
    pxcRom[6890] <= 10'b0000000000;
    pxcRom[6891] <= 10'b0000000000;
    pxcRom[6892] <= 10'b0000000000;
    pxcRom[6893] <= 10'b0000000011;
    pxcRom[6894] <= 10'b0000001010;
    pxcRom[6895] <= 10'b0000010101;
    pxcRom[6896] <= 10'b0000100110;
    pxcRom[6897] <= 10'b0000111011;
    pxcRom[6898] <= 10'b0001010110;
    pxcRom[6899] <= 10'b0001101100;
    pxcRom[6900] <= 10'b0001110100;
    pxcRom[6901] <= 10'b0001110100;
    pxcRom[6902] <= 10'b0001101011;
    pxcRom[6903] <= 10'b0001010111;
    pxcRom[6904] <= 10'b0001000000;
    pxcRom[6905] <= 10'b0000101011;
    pxcRom[6906] <= 10'b0000011011;
    pxcRom[6907] <= 10'b0000001111;
    pxcRom[6908] <= 10'b0000001000;
    pxcRom[6909] <= 10'b0000000011;
    pxcRom[6910] <= 10'b0000000001;
    pxcRom[6911] <= 10'b0000000000;
    pxcRom[6912] <= 10'b0000000000;
    pxcRom[6913] <= 10'b0000000000;
    pxcRom[6914] <= 10'b0000000000;
    pxcRom[6915] <= 10'b0000000000;
    pxcRom[6916] <= 10'b0000000000;
    pxcRom[6917] <= 10'b0000000000;
    pxcRom[6918] <= 10'b0000000000;
    pxcRom[6919] <= 10'b0000000000;
    pxcRom[6920] <= 10'b0000000000;
    pxcRom[6921] <= 10'b0000000010;
    pxcRom[6922] <= 10'b0000000111;
    pxcRom[6923] <= 10'b0000001111;
    pxcRom[6924] <= 10'b0000011100;
    pxcRom[6925] <= 10'b0000101101;
    pxcRom[6926] <= 10'b0001000100;
    pxcRom[6927] <= 10'b0001100011;
    pxcRom[6928] <= 10'b0001111000;
    pxcRom[6929] <= 10'b0001110110;
    pxcRom[6930] <= 10'b0001100010;
    pxcRom[6931] <= 10'b0001000110;
    pxcRom[6932] <= 10'b0000101111;
    pxcRom[6933] <= 10'b0000011101;
    pxcRom[6934] <= 10'b0000010000;
    pxcRom[6935] <= 10'b0000001000;
    pxcRom[6936] <= 10'b0000000100;
    pxcRom[6937] <= 10'b0000000001;
    pxcRom[6938] <= 10'b0000000000;
    pxcRom[6939] <= 10'b0000000000;
    pxcRom[6940] <= 10'b0000000000;
    pxcRom[6941] <= 10'b0000000000;
    pxcRom[6942] <= 10'b0000000000;
    pxcRom[6943] <= 10'b0000000000;
    pxcRom[6944] <= 10'b0000000000;
    pxcRom[6945] <= 10'b0000000000;
    pxcRom[6946] <= 10'b0000000000;
    pxcRom[6947] <= 10'b0000000000;
    pxcRom[6948] <= 10'b0000000000;
    pxcRom[6949] <= 10'b0000000000;
    pxcRom[6950] <= 10'b0000000010;
    pxcRom[6951] <= 10'b0000000110;
    pxcRom[6952] <= 10'b0000001100;
    pxcRom[6953] <= 10'b0000010101;
    pxcRom[6954] <= 10'b0000011111;
    pxcRom[6955] <= 10'b0000101001;
    pxcRom[6956] <= 10'b0000101111;
    pxcRom[6957] <= 10'b0000101110;
    pxcRom[6958] <= 10'b0000100110;
    pxcRom[6959] <= 10'b0000011101;
    pxcRom[6960] <= 10'b0000010011;
    pxcRom[6961] <= 10'b0000001011;
    pxcRom[6962] <= 10'b0000000110;
    pxcRom[6963] <= 10'b0000000011;
    pxcRom[6964] <= 10'b0000000001;
    pxcRom[6965] <= 10'b0000000000;
    pxcRom[6966] <= 10'b0000000000;
    pxcRom[6967] <= 10'b0000000000;
    pxcRom[6968] <= 10'b0000000000;
    pxcRom[6969] <= 10'b0000000000;
    pxcRom[6970] <= 10'b0000000000;
    pxcRom[6971] <= 10'b0000000000;
    pxcRom[6972] <= 10'b0000000000;
    pxcRom[6973] <= 10'b0000000000;
    pxcRom[6974] <= 10'b0000000000;
    pxcRom[6975] <= 10'b0000000000;
    pxcRom[6976] <= 10'b0000000000;
    pxcRom[6977] <= 10'b0000000000;
    pxcRom[6978] <= 10'b0000000000;
    pxcRom[6979] <= 10'b0000000000;
    pxcRom[6980] <= 10'b0000000001;
    pxcRom[6981] <= 10'b0000000001;
    pxcRom[6982] <= 10'b0000000010;
    pxcRom[6983] <= 10'b0000000010;
    pxcRom[6984] <= 10'b0000000011;
    pxcRom[6985] <= 10'b0000000011;
    pxcRom[6986] <= 10'b0000000011;
    pxcRom[6987] <= 10'b0000000010;
    pxcRom[6988] <= 10'b0000000001;
    pxcRom[6989] <= 10'b0000000001;
    pxcRom[6990] <= 10'b0000000000;
    pxcRom[6991] <= 10'b0000000000;
    pxcRom[6992] <= 10'b0000000000;
    pxcRom[6993] <= 10'b0000000000;
    pxcRom[6994] <= 10'b0000000000;
    pxcRom[6995] <= 10'b0000000000;
    pxcRom[6996] <= 10'b0000000000;
    pxcRom[6997] <= 10'b0000000000;
    pxcRom[6998] <= 10'b0000000000;
    pxcRom[6999] <= 10'b0000000000;
    pxcRom[7000] <= 10'b0000000000;
    pxcRom[7001] <= 10'b0000000000;
    pxcRom[7002] <= 10'b0000000000;
    pxcRom[7003] <= 10'b0000000000;
    pxcRom[7004] <= 10'b0000000000;
    pxcRom[7005] <= 10'b0000000000;
    pxcRom[7006] <= 10'b0000000000;
    pxcRom[7007] <= 10'b0000000000;
    pxcRom[7008] <= 10'b0000000000;
    pxcRom[7009] <= 10'b0000000000;
    pxcRom[7010] <= 10'b0000000000;
    pxcRom[7011] <= 10'b0000000000;
    pxcRom[7012] <= 10'b0000000000;
    pxcRom[7013] <= 10'b0000000000;
    pxcRom[7014] <= 10'b0000000000;
    pxcRom[7015] <= 10'b0000000000;
    pxcRom[7016] <= 10'b0000000000;
    pxcRom[7017] <= 10'b0000000000;
    pxcRom[7018] <= 10'b0000000000;
    pxcRom[7019] <= 10'b0000000000;
    pxcRom[7020] <= 10'b0000000000;
    pxcRom[7021] <= 10'b0000000000;
    pxcRom[7022] <= 10'b0000000000;
    pxcRom[7023] <= 10'b0000000000;
    pxcRom[7024] <= 10'b0000000000;
    pxcRom[7025] <= 10'b0000000000;
    pxcRom[7026] <= 10'b0000000000;
    pxcRom[7027] <= 10'b0000000000;
    pxcRom[7028] <= 10'b0000000000;
    pxcRom[7029] <= 10'b0000000000;
    pxcRom[7030] <= 10'b0000000000;
    pxcRom[7031] <= 10'b0000000000;
    pxcRom[7032] <= 10'b0000000000;
    pxcRom[7033] <= 10'b0000000000;
    pxcRom[7034] <= 10'b0000000000;
    pxcRom[7035] <= 10'b0000000000;
    pxcRom[7036] <= 10'b0000000000;
    pxcRom[7037] <= 10'b0000000000;
    pxcRom[7038] <= 10'b0000000000;
    pxcRom[7039] <= 10'b0000000000;
    pxcRom[7040] <= 10'b0000000000;
    pxcRom[7041] <= 10'b0000000000;
    pxcRom[7042] <= 10'b0000000000;
    pxcRom[7043] <= 10'b0000000000;
    pxcRom[7044] <= 10'b0000000000;
    pxcRom[7045] <= 10'b0000000000;
    pxcRom[7046] <= 10'b0000000000;
    pxcRom[7047] <= 10'b0000000000;
    pxcRom[7048] <= 10'b0000000000;
    pxcRom[7049] <= 10'b0000000000;
    pxcRom[7050] <= 10'b0000000000;
    pxcRom[7051] <= 10'b0000000000;
    pxcRom[7052] <= 10'b0000000000;
    pxcRom[7053] <= 10'b0000000000;
    pxcRom[7054] <= 10'b0000000000;
    pxcRom[7055] <= 10'b0000000000;
    pxcRom[7056] <= 10'b0000000000;
    pxcRom[7057] <= 10'b0000000000;
    pxcRom[7058] <= 10'b0000000000;
    pxcRom[7059] <= 10'b0000000000;
    pxcRom[7060] <= 10'b0000000000;
    pxcRom[7061] <= 10'b0000000000;
    pxcRom[7062] <= 10'b0000000000;
    pxcRom[7063] <= 10'b0000000000;
    pxcRom[7064] <= 10'b0000000000;
    pxcRom[7065] <= 10'b0000000000;
    pxcRom[7066] <= 10'b0000000000;
    pxcRom[7067] <= 10'b0000000000;
    pxcRom[7068] <= 10'b0000000000;
    pxcRom[7069] <= 10'b0000000000;
    pxcRom[7070] <= 10'b0000000000;
    pxcRom[7071] <= 10'b0000000000;
    pxcRom[7072] <= 10'b0000000000;
    pxcRom[7073] <= 10'b0000000000;
    pxcRom[7074] <= 10'b0000000000;
    pxcRom[7075] <= 10'b0000000000;
    pxcRom[7076] <= 10'b0000000000;
    pxcRom[7077] <= 10'b0000000000;
    pxcRom[7078] <= 10'b0000000000;
    pxcRom[7079] <= 10'b0000000000;
    pxcRom[7080] <= 10'b0000000000;
    pxcRom[7081] <= 10'b0000000000;
    pxcRom[7082] <= 10'b0000000000;
    pxcRom[7083] <= 10'b0000000000;
    pxcRom[7084] <= 10'b0000000000;
    pxcRom[7085] <= 10'b0000000000;
    pxcRom[7086] <= 10'b0000000000;
    pxcRom[7087] <= 10'b0000000000;
    pxcRom[7088] <= 10'b0000000000;
    pxcRom[7089] <= 10'b0000000000;
    pxcRom[7090] <= 10'b0000000000;
    pxcRom[7091] <= 10'b0000000000;
    pxcRom[7092] <= 10'b0000000000;
    pxcRom[7093] <= 10'b0000000000;
    pxcRom[7094] <= 10'b0000000000;
    pxcRom[7095] <= 10'b0000000000;
    pxcRom[7096] <= 10'b0000000000;
    pxcRom[7097] <= 10'b0000000000;
    pxcRom[7098] <= 10'b0000000000;
    pxcRom[7099] <= 10'b0000000000;
    pxcRom[7100] <= 10'b0000000000;
    pxcRom[7101] <= 10'b0000000000;
    pxcRom[7102] <= 10'b0000000000;
    pxcRom[7103] <= 10'b0000000000;
    pxcRom[7104] <= 10'b0000000000;
    pxcRom[7105] <= 10'b0000000000;
    pxcRom[7106] <= 10'b0000000000;
    pxcRom[7107] <= 10'b0000000000;
    pxcRom[7108] <= 10'b0000000000;
    pxcRom[7109] <= 10'b0000000000;
    pxcRom[7110] <= 10'b0000000000;
    pxcRom[7111] <= 10'b0000000000;
    pxcRom[7112] <= 10'b0000000000;
    pxcRom[7113] <= 10'b0000000000;
    pxcRom[7114] <= 10'b0000000000;
    pxcRom[7115] <= 10'b0000000000;
    pxcRom[7116] <= 10'b0000000000;
    pxcRom[7117] <= 10'b0000000000;
    pxcRom[7118] <= 10'b0000000000;
    pxcRom[7119] <= 10'b0000000000;
    pxcRom[7120] <= 10'b0000000000;
    pxcRom[7121] <= 10'b0000000000;
    pxcRom[7122] <= 10'b0000000000;
    pxcRom[7123] <= 10'b0000000000;
    pxcRom[7124] <= 10'b0000000000;
    pxcRom[7125] <= 10'b0000000000;
    pxcRom[7126] <= 10'b0000000000;
    pxcRom[7127] <= 10'b0000000000;
    pxcRom[7128] <= 10'b0000000000;
    pxcRom[7129] <= 10'b0000000000;
    pxcRom[7130] <= 10'b0000000000;
    pxcRom[7131] <= 10'b0000000000;
    pxcRom[7132] <= 10'b0000000000;
    pxcRom[7133] <= 10'b0000000000;
    pxcRom[7134] <= 10'b0000000000;
    pxcRom[7135] <= 10'b0000000000;
    pxcRom[7136] <= 10'b0000000000;
    pxcRom[7137] <= 10'b0000000000;
    pxcRom[7138] <= 10'b0000000000;
    pxcRom[7139] <= 10'b0000000000;
    pxcRom[7140] <= 10'b0000000000;
    pxcRom[7141] <= 10'b0000000000;
    pxcRom[7142] <= 10'b0000000000;
    pxcRom[7143] <= 10'b0000000000;
    pxcRom[7144] <= 10'b0000000000;
    pxcRom[7145] <= 10'b0000000000;
    pxcRom[7146] <= 10'b0000000000;
    pxcRom[7147] <= 10'b0000000000;
    pxcRom[7148] <= 10'b0000000000;
    pxcRom[7149] <= 10'b0000000000;
    pxcRom[7150] <= 10'b0000000000;
    pxcRom[7151] <= 10'b0000000000;
    pxcRom[7152] <= 10'b0000000000;
    pxcRom[7153] <= 10'b0000000000;
    pxcRom[7154] <= 10'b0000000000;
    pxcRom[7155] <= 10'b0000000000;
    pxcRom[7156] <= 10'b0000000000;
    pxcRom[7157] <= 10'b0000000000;
    pxcRom[7158] <= 10'b0000000000;
    pxcRom[7159] <= 10'b0000000000;
    pxcRom[7160] <= 10'b0000000000;
    pxcRom[7161] <= 10'b0000000000;
    pxcRom[7162] <= 10'b0000000000;
    pxcRom[7163] <= 10'b0000000000;
    pxcRom[7164] <= 10'b0000000000;
    pxcRom[7165] <= 10'b0000000000;
    pxcRom[7166] <= 10'b0000000000;
    pxcRom[7167] <= 10'b0000000000;
    pxcRom[7168] <= 10'b0000000000;
    pxcRom[7169] <= 10'b0000000000;
    pxcRom[7170] <= 10'b0000000000;
    pxcRom[7171] <= 10'b0000000000;
    pxcRom[7172] <= 10'b0000000000;
    pxcRom[7173] <= 10'b0000000000;
    pxcRom[7174] <= 10'b0000000000;
    pxcRom[7175] <= 10'b0000000000;
    pxcRom[7176] <= 10'b0000000000;
    pxcRom[7177] <= 10'b0000000000;
    pxcRom[7178] <= 10'b0000000000;
    pxcRom[7179] <= 10'b0000000000;
    pxcRom[7180] <= 10'b0000000000;
    pxcRom[7181] <= 10'b0000000000;
    pxcRom[7182] <= 10'b0000000000;
    pxcRom[7183] <= 10'b0000000000;
    pxcRom[7184] <= 10'b0000000000;
    pxcRom[7185] <= 10'b0000000000;
    pxcRom[7186] <= 10'b0000000000;
    pxcRom[7187] <= 10'b0000000000;
    pxcRom[7188] <= 10'b0000000000;
    pxcRom[7189] <= 10'b0000000000;
    pxcRom[7190] <= 10'b0000000000;
    pxcRom[7191] <= 10'b0000000000;
    pxcRom[7192] <= 10'b0000000000;
    pxcRom[7193] <= 10'b0000000000;
    pxcRom[7194] <= 10'b0000000000;
    pxcRom[7195] <= 10'b0000000000;
    pxcRom[7196] <= 10'b0000000000;
    pxcRom[7197] <= 10'b0000000000;
    pxcRom[7198] <= 10'b0000000000;
    pxcRom[7199] <= 10'b0000000000;
    pxcRom[7200] <= 10'b0000000000;
    pxcRom[7201] <= 10'b0000000000;
    pxcRom[7202] <= 10'b0000000000;
    pxcRom[7203] <= 10'b0000000000;
    pxcRom[7204] <= 10'b0000000000;
    pxcRom[7205] <= 10'b0000000000;
    pxcRom[7206] <= 10'b0000000000;
    pxcRom[7207] <= 10'b0000000001;
    pxcRom[7208] <= 10'b0000000010;
    pxcRom[7209] <= 10'b0000000011;
    pxcRom[7210] <= 10'b0000000011;
    pxcRom[7211] <= 10'b0000000100;
    pxcRom[7212] <= 10'b0000000011;
    pxcRom[7213] <= 10'b0000000010;
    pxcRom[7214] <= 10'b0000000001;
    pxcRom[7215] <= 10'b0000000001;
    pxcRom[7216] <= 10'b0000000000;
    pxcRom[7217] <= 10'b0000000000;
    pxcRom[7218] <= 10'b0000000000;
    pxcRom[7219] <= 10'b0000000000;
    pxcRom[7220] <= 10'b0000000000;
    pxcRom[7221] <= 10'b0000000000;
    pxcRom[7222] <= 10'b0000000000;
    pxcRom[7223] <= 10'b0000000000;
    pxcRom[7224] <= 10'b0000000000;
    pxcRom[7225] <= 10'b0000000000;
    pxcRom[7226] <= 10'b0000000000;
    pxcRom[7227] <= 10'b0000000000;
    pxcRom[7228] <= 10'b0000000000;
    pxcRom[7229] <= 10'b0000000000;
    pxcRom[7230] <= 10'b0000000000;
    pxcRom[7231] <= 10'b0000000000;
    pxcRom[7232] <= 10'b0000000001;
    pxcRom[7233] <= 10'b0000000011;
    pxcRom[7234] <= 10'b0000000110;
    pxcRom[7235] <= 10'b0000001101;
    pxcRom[7236] <= 10'b0000011000;
    pxcRom[7237] <= 10'b0000100100;
    pxcRom[7238] <= 10'b0000110000;
    pxcRom[7239] <= 10'b0000110111;
    pxcRom[7240] <= 10'b0000110010;
    pxcRom[7241] <= 10'b0000100111;
    pxcRom[7242] <= 10'b0000011010;
    pxcRom[7243] <= 10'b0000001111;
    pxcRom[7244] <= 10'b0000000111;
    pxcRom[7245] <= 10'b0000000011;
    pxcRom[7246] <= 10'b0000000001;
    pxcRom[7247] <= 10'b0000000000;
    pxcRom[7248] <= 10'b0000000000;
    pxcRom[7249] <= 10'b0000000000;
    pxcRom[7250] <= 10'b0000000000;
    pxcRom[7251] <= 10'b0000000000;
    pxcRom[7252] <= 10'b0000000000;
    pxcRom[7253] <= 10'b0000000000;
    pxcRom[7254] <= 10'b0000000000;
    pxcRom[7255] <= 10'b0000000000;
    pxcRom[7256] <= 10'b0000000000;
    pxcRom[7257] <= 10'b0000000000;
    pxcRom[7258] <= 10'b0000000000;
    pxcRom[7259] <= 10'b0000000010;
    pxcRom[7260] <= 10'b0000000101;
    pxcRom[7261] <= 10'b0000001011;
    pxcRom[7262] <= 10'b0000011000;
    pxcRom[7263] <= 10'b0000101100;
    pxcRom[7264] <= 10'b0001001011;
    pxcRom[7265] <= 10'b0001110100;
    pxcRom[7266] <= 10'b0010010110;
    pxcRom[7267] <= 10'b0010100010;
    pxcRom[7268] <= 10'b0010000110;
    pxcRom[7269] <= 10'b0001011110;
    pxcRom[7270] <= 10'b0000111100;
    pxcRom[7271] <= 10'b0000100010;
    pxcRom[7272] <= 10'b0000010001;
    pxcRom[7273] <= 10'b0000001000;
    pxcRom[7274] <= 10'b0000000011;
    pxcRom[7275] <= 10'b0000000000;
    pxcRom[7276] <= 10'b0000000000;
    pxcRom[7277] <= 10'b0000000000;
    pxcRom[7278] <= 10'b0000000000;
    pxcRom[7279] <= 10'b0000000000;
    pxcRom[7280] <= 10'b0000000000;
    pxcRom[7281] <= 10'b0000000000;
    pxcRom[7282] <= 10'b0000000000;
    pxcRom[7283] <= 10'b0000000000;
    pxcRom[7284] <= 10'b0000000000;
    pxcRom[7285] <= 10'b0000000000;
    pxcRom[7286] <= 10'b0000000010;
    pxcRom[7287] <= 10'b0000000101;
    pxcRom[7288] <= 10'b0000001101;
    pxcRom[7289] <= 10'b0000011100;
    pxcRom[7290] <= 10'b0000110110;
    pxcRom[7291] <= 10'b0001011101;
    pxcRom[7292] <= 10'b0010000001;
    pxcRom[7293] <= 10'b0010001000;
    pxcRom[7294] <= 10'b0001111101;
    pxcRom[7295] <= 10'b0001110101;
    pxcRom[7296] <= 10'b0001110001;
    pxcRom[7297] <= 10'b0001100110;
    pxcRom[7298] <= 10'b0001001110;
    pxcRom[7299] <= 10'b0000101111;
    pxcRom[7300] <= 10'b0000011010;
    pxcRom[7301] <= 10'b0000001100;
    pxcRom[7302] <= 10'b0000000101;
    pxcRom[7303] <= 10'b0000000001;
    pxcRom[7304] <= 10'b0000000000;
    pxcRom[7305] <= 10'b0000000000;
    pxcRom[7306] <= 10'b0000000000;
    pxcRom[7307] <= 10'b0000000000;
    pxcRom[7308] <= 10'b0000000000;
    pxcRom[7309] <= 10'b0000000000;
    pxcRom[7310] <= 10'b0000000000;
    pxcRom[7311] <= 10'b0000000000;
    pxcRom[7312] <= 10'b0000000000;
    pxcRom[7313] <= 10'b0000000001;
    pxcRom[7314] <= 10'b0000000100;
    pxcRom[7315] <= 10'b0000001011;
    pxcRom[7316] <= 10'b0000011010;
    pxcRom[7317] <= 10'b0000110100;
    pxcRom[7318] <= 10'b0001011001;
    pxcRom[7319] <= 10'b0001110000;
    pxcRom[7320] <= 10'b0001100000;
    pxcRom[7321] <= 10'b0001000101;
    pxcRom[7322] <= 10'b0000110100;
    pxcRom[7323] <= 10'b0000110000;
    pxcRom[7324] <= 10'b0000111011;
    pxcRom[7325] <= 10'b0001001011;
    pxcRom[7326] <= 10'b0001001101;
    pxcRom[7327] <= 10'b0000111001;
    pxcRom[7328] <= 10'b0000011111;
    pxcRom[7329] <= 10'b0000001111;
    pxcRom[7330] <= 10'b0000000110;
    pxcRom[7331] <= 10'b0000000001;
    pxcRom[7332] <= 10'b0000000000;
    pxcRom[7333] <= 10'b0000000000;
    pxcRom[7334] <= 10'b0000000000;
    pxcRom[7335] <= 10'b0000000000;
    pxcRom[7336] <= 10'b0000000000;
    pxcRom[7337] <= 10'b0000000000;
    pxcRom[7338] <= 10'b0000000000;
    pxcRom[7339] <= 10'b0000000000;
    pxcRom[7340] <= 10'b0000000001;
    pxcRom[7341] <= 10'b0000000011;
    pxcRom[7342] <= 10'b0000001000;
    pxcRom[7343] <= 10'b0000010100;
    pxcRom[7344] <= 10'b0000101010;
    pxcRom[7345] <= 10'b0001001101;
    pxcRom[7346] <= 10'b0001100100;
    pxcRom[7347] <= 10'b0001010001;
    pxcRom[7348] <= 10'b0000110001;
    pxcRom[7349] <= 10'b0000011011;
    pxcRom[7350] <= 10'b0000010011;
    pxcRom[7351] <= 10'b0000011000;
    pxcRom[7352] <= 10'b0000101010;
    pxcRom[7353] <= 10'b0001000111;
    pxcRom[7354] <= 10'b0001010101;
    pxcRom[7355] <= 10'b0001000001;
    pxcRom[7356] <= 10'b0000100011;
    pxcRom[7357] <= 10'b0000010000;
    pxcRom[7358] <= 10'b0000000110;
    pxcRom[7359] <= 10'b0000000001;
    pxcRom[7360] <= 10'b0000000000;
    pxcRom[7361] <= 10'b0000000000;
    pxcRom[7362] <= 10'b0000000000;
    pxcRom[7363] <= 10'b0000000000;
    pxcRom[7364] <= 10'b0000000000;
    pxcRom[7365] <= 10'b0000000000;
    pxcRom[7366] <= 10'b0000000000;
    pxcRom[7367] <= 10'b0000000000;
    pxcRom[7368] <= 10'b0000000001;
    pxcRom[7369] <= 10'b0000000101;
    pxcRom[7370] <= 10'b0000001100;
    pxcRom[7371] <= 10'b0000011101;
    pxcRom[7372] <= 10'b0000111010;
    pxcRom[7373] <= 10'b0001011010;
    pxcRom[7374] <= 10'b0001010100;
    pxcRom[7375] <= 10'b0000110010;
    pxcRom[7376] <= 10'b0000011000;
    pxcRom[7377] <= 10'b0000001100;
    pxcRom[7378] <= 10'b0000001100;
    pxcRom[7379] <= 10'b0000011010;
    pxcRom[7380] <= 10'b0000110100;
    pxcRom[7381] <= 10'b0001011010;
    pxcRom[7382] <= 10'b0001101000;
    pxcRom[7383] <= 10'b0001000110;
    pxcRom[7384] <= 10'b0000100011;
    pxcRom[7385] <= 10'b0000001110;
    pxcRom[7386] <= 10'b0000000101;
    pxcRom[7387] <= 10'b0000000001;
    pxcRom[7388] <= 10'b0000000000;
    pxcRom[7389] <= 10'b0000000000;
    pxcRom[7390] <= 10'b0000000000;
    pxcRom[7391] <= 10'b0000000000;
    pxcRom[7392] <= 10'b0000000000;
    pxcRom[7393] <= 10'b0000000000;
    pxcRom[7394] <= 10'b0000000000;
    pxcRom[7395] <= 10'b0000000000;
    pxcRom[7396] <= 10'b0000000010;
    pxcRom[7397] <= 10'b0000000110;
    pxcRom[7398] <= 10'b0000001111;
    pxcRom[7399] <= 10'b0000100100;
    pxcRom[7400] <= 10'b0001000011;
    pxcRom[7401] <= 10'b0001011000;
    pxcRom[7402] <= 10'b0001000011;
    pxcRom[7403] <= 10'b0000100011;
    pxcRom[7404] <= 10'b0000010001;
    pxcRom[7405] <= 10'b0000001111;
    pxcRom[7406] <= 10'b0000011000;
    pxcRom[7407] <= 10'b0000101101;
    pxcRom[7408] <= 10'b0001010010;
    pxcRom[7409] <= 10'b0001111110;
    pxcRom[7410] <= 10'b0001110100;
    pxcRom[7411] <= 10'b0001000001;
    pxcRom[7412] <= 10'b0000011110;
    pxcRom[7413] <= 10'b0000001011;
    pxcRom[7414] <= 10'b0000000100;
    pxcRom[7415] <= 10'b0000000001;
    pxcRom[7416] <= 10'b0000000000;
    pxcRom[7417] <= 10'b0000000000;
    pxcRom[7418] <= 10'b0000000000;
    pxcRom[7419] <= 10'b0000000000;
    pxcRom[7420] <= 10'b0000000000;
    pxcRom[7421] <= 10'b0000000000;
    pxcRom[7422] <= 10'b0000000000;
    pxcRom[7423] <= 10'b0000000000;
    pxcRom[7424] <= 10'b0000000010;
    pxcRom[7425] <= 10'b0000000111;
    pxcRom[7426] <= 10'b0000010001;
    pxcRom[7427] <= 10'b0000100110;
    pxcRom[7428] <= 10'b0001000100;
    pxcRom[7429] <= 10'b0001010010;
    pxcRom[7430] <= 10'b0000111110;
    pxcRom[7431] <= 10'b0000100110;
    pxcRom[7432] <= 10'b0000011110;
    pxcRom[7433] <= 10'b0000100011;
    pxcRom[7434] <= 10'b0000110011;
    pxcRom[7435] <= 10'b0001010000;
    pxcRom[7436] <= 10'b0001111101;
    pxcRom[7437] <= 10'b0010100000;
    pxcRom[7438] <= 10'b0001101110;
    pxcRom[7439] <= 10'b0000110110;
    pxcRom[7440] <= 10'b0000010110;
    pxcRom[7441] <= 10'b0000001000;
    pxcRom[7442] <= 10'b0000000010;
    pxcRom[7443] <= 10'b0000000000;
    pxcRom[7444] <= 10'b0000000000;
    pxcRom[7445] <= 10'b0000000000;
    pxcRom[7446] <= 10'b0000000000;
    pxcRom[7447] <= 10'b0000000000;
    pxcRom[7448] <= 10'b0000000000;
    pxcRom[7449] <= 10'b0000000000;
    pxcRom[7450] <= 10'b0000000000;
    pxcRom[7451] <= 10'b0000000000;
    pxcRom[7452] <= 10'b0000000010;
    pxcRom[7453] <= 10'b0000000111;
    pxcRom[7454] <= 10'b0000010000;
    pxcRom[7455] <= 10'b0000100011;
    pxcRom[7456] <= 10'b0000111110;
    pxcRom[7457] <= 10'b0001001111;
    pxcRom[7458] <= 10'b0001000111;
    pxcRom[7459] <= 10'b0000111011;
    pxcRom[7460] <= 10'b0000111010;
    pxcRom[7461] <= 10'b0001000011;
    pxcRom[7462] <= 10'b0001010100;
    pxcRom[7463] <= 10'b0001101110;
    pxcRom[7464] <= 10'b0010011110;
    pxcRom[7465] <= 10'b0010101000;
    pxcRom[7466] <= 10'b0001011100;
    pxcRom[7467] <= 10'b0000100111;
    pxcRom[7468] <= 10'b0000001110;
    pxcRom[7469] <= 10'b0000000101;
    pxcRom[7470] <= 10'b0000000001;
    pxcRom[7471] <= 10'b0000000000;
    pxcRom[7472] <= 10'b0000000000;
    pxcRom[7473] <= 10'b0000000000;
    pxcRom[7474] <= 10'b0000000000;
    pxcRom[7475] <= 10'b0000000000;
    pxcRom[7476] <= 10'b0000000000;
    pxcRom[7477] <= 10'b0000000000;
    pxcRom[7478] <= 10'b0000000000;
    pxcRom[7479] <= 10'b0000000000;
    pxcRom[7480] <= 10'b0000000001;
    pxcRom[7481] <= 10'b0000000101;
    pxcRom[7482] <= 10'b0000001101;
    pxcRom[7483] <= 10'b0000011011;
    pxcRom[7484] <= 10'b0000110001;
    pxcRom[7485] <= 10'b0001000100;
    pxcRom[7486] <= 10'b0001001100;
    pxcRom[7487] <= 10'b0001001011;
    pxcRom[7488] <= 10'b0001001100;
    pxcRom[7489] <= 10'b0001001111;
    pxcRom[7490] <= 10'b0001010111;
    pxcRom[7491] <= 10'b0001110011;
    pxcRom[7492] <= 10'b0010100000;
    pxcRom[7493] <= 10'b0010010000;
    pxcRom[7494] <= 10'b0001000110;
    pxcRom[7495] <= 10'b0000011011;
    pxcRom[7496] <= 10'b0000001010;
    pxcRom[7497] <= 10'b0000000011;
    pxcRom[7498] <= 10'b0000000001;
    pxcRom[7499] <= 10'b0000000000;
    pxcRom[7500] <= 10'b0000000000;
    pxcRom[7501] <= 10'b0000000000;
    pxcRom[7502] <= 10'b0000000000;
    pxcRom[7503] <= 10'b0000000000;
    pxcRom[7504] <= 10'b0000000000;
    pxcRom[7505] <= 10'b0000000000;
    pxcRom[7506] <= 10'b0000000000;
    pxcRom[7507] <= 10'b0000000000;
    pxcRom[7508] <= 10'b0000000001;
    pxcRom[7509] <= 10'b0000000011;
    pxcRom[7510] <= 10'b0000001000;
    pxcRom[7511] <= 10'b0000010010;
    pxcRom[7512] <= 10'b0000100000;
    pxcRom[7513] <= 10'b0000101111;
    pxcRom[7514] <= 10'b0000111001;
    pxcRom[7515] <= 10'b0000111101;
    pxcRom[7516] <= 10'b0000111101;
    pxcRom[7517] <= 10'b0000111011;
    pxcRom[7518] <= 10'b0001000111;
    pxcRom[7519] <= 10'b0001100110;
    pxcRom[7520] <= 10'b0010001101;
    pxcRom[7521] <= 10'b0001101101;
    pxcRom[7522] <= 10'b0000110010;
    pxcRom[7523] <= 10'b0000010011;
    pxcRom[7524] <= 10'b0000000111;
    pxcRom[7525] <= 10'b0000000010;
    pxcRom[7526] <= 10'b0000000001;
    pxcRom[7527] <= 10'b0000000000;
    pxcRom[7528] <= 10'b0000000000;
    pxcRom[7529] <= 10'b0000000000;
    pxcRom[7530] <= 10'b0000000000;
    pxcRom[7531] <= 10'b0000000000;
    pxcRom[7532] <= 10'b0000000000;
    pxcRom[7533] <= 10'b0000000000;
    pxcRom[7534] <= 10'b0000000000;
    pxcRom[7535] <= 10'b0000000000;
    pxcRom[7536] <= 10'b0000000000;
    pxcRom[7537] <= 10'b0000000010;
    pxcRom[7538] <= 10'b0000000100;
    pxcRom[7539] <= 10'b0000001001;
    pxcRom[7540] <= 10'b0000010000;
    pxcRom[7541] <= 10'b0000011000;
    pxcRom[7542] <= 10'b0000011110;
    pxcRom[7543] <= 10'b0000100000;
    pxcRom[7544] <= 10'b0000100001;
    pxcRom[7545] <= 10'b0000100110;
    pxcRom[7546] <= 10'b0000111011;
    pxcRom[7547] <= 10'b0001011101;
    pxcRom[7548] <= 10'b0001110010;
    pxcRom[7549] <= 10'b0001001111;
    pxcRom[7550] <= 10'b0000100100;
    pxcRom[7551] <= 10'b0000001111;
    pxcRom[7552] <= 10'b0000000110;
    pxcRom[7553] <= 10'b0000000010;
    pxcRom[7554] <= 10'b0000000000;
    pxcRom[7555] <= 10'b0000000000;
    pxcRom[7556] <= 10'b0000000000;
    pxcRom[7557] <= 10'b0000000000;
    pxcRom[7558] <= 10'b0000000000;
    pxcRom[7559] <= 10'b0000000000;
    pxcRom[7560] <= 10'b0000000000;
    pxcRom[7561] <= 10'b0000000000;
    pxcRom[7562] <= 10'b0000000000;
    pxcRom[7563] <= 10'b0000000000;
    pxcRom[7564] <= 10'b0000000000;
    pxcRom[7565] <= 10'b0000000000;
    pxcRom[7566] <= 10'b0000000010;
    pxcRom[7567] <= 10'b0000000100;
    pxcRom[7568] <= 10'b0000000111;
    pxcRom[7569] <= 10'b0000001010;
    pxcRom[7570] <= 10'b0000001101;
    pxcRom[7571] <= 10'b0000001111;
    pxcRom[7572] <= 10'b0000010011;
    pxcRom[7573] <= 10'b0000011110;
    pxcRom[7574] <= 10'b0000110110;
    pxcRom[7575] <= 10'b0001010010;
    pxcRom[7576] <= 10'b0001010111;
    pxcRom[7577] <= 10'b0000111000;
    pxcRom[7578] <= 10'b0000011100;
    pxcRom[7579] <= 10'b0000001100;
    pxcRom[7580] <= 10'b0000000101;
    pxcRom[7581] <= 10'b0000000010;
    pxcRom[7582] <= 10'b0000000001;
    pxcRom[7583] <= 10'b0000000000;
    pxcRom[7584] <= 10'b0000000000;
    pxcRom[7585] <= 10'b0000000000;
    pxcRom[7586] <= 10'b0000000000;
    pxcRom[7587] <= 10'b0000000000;
    pxcRom[7588] <= 10'b0000000000;
    pxcRom[7589] <= 10'b0000000000;
    pxcRom[7590] <= 10'b0000000000;
    pxcRom[7591] <= 10'b0000000000;
    pxcRom[7592] <= 10'b0000000000;
    pxcRom[7593] <= 10'b0000000000;
    pxcRom[7594] <= 10'b0000000000;
    pxcRom[7595] <= 10'b0000000001;
    pxcRom[7596] <= 10'b0000000010;
    pxcRom[7597] <= 10'b0000000011;
    pxcRom[7598] <= 10'b0000000101;
    pxcRom[7599] <= 10'b0000001000;
    pxcRom[7600] <= 10'b0000010000;
    pxcRom[7601] <= 10'b0000011111;
    pxcRom[7602] <= 10'b0000110101;
    pxcRom[7603] <= 10'b0001000111;
    pxcRom[7604] <= 10'b0001000011;
    pxcRom[7605] <= 10'b0000101010;
    pxcRom[7606] <= 10'b0000010111;
    pxcRom[7607] <= 10'b0000001011;
    pxcRom[7608] <= 10'b0000000101;
    pxcRom[7609] <= 10'b0000000010;
    pxcRom[7610] <= 10'b0000000001;
    pxcRom[7611] <= 10'b0000000000;
    pxcRom[7612] <= 10'b0000000000;
    pxcRom[7613] <= 10'b0000000000;
    pxcRom[7614] <= 10'b0000000000;
    pxcRom[7615] <= 10'b0000000000;
    pxcRom[7616] <= 10'b0000000000;
    pxcRom[7617] <= 10'b0000000000;
    pxcRom[7618] <= 10'b0000000000;
    pxcRom[7619] <= 10'b0000000000;
    pxcRom[7620] <= 10'b0000000000;
    pxcRom[7621] <= 10'b0000000000;
    pxcRom[7622] <= 10'b0000000000;
    pxcRom[7623] <= 10'b0000000000;
    pxcRom[7624] <= 10'b0000000001;
    pxcRom[7625] <= 10'b0000000010;
    pxcRom[7626] <= 10'b0000000100;
    pxcRom[7627] <= 10'b0000001001;
    pxcRom[7628] <= 10'b0000010100;
    pxcRom[7629] <= 10'b0000100100;
    pxcRom[7630] <= 10'b0000110100;
    pxcRom[7631] <= 10'b0000111100;
    pxcRom[7632] <= 10'b0000110010;
    pxcRom[7633] <= 10'b0000100010;
    pxcRom[7634] <= 10'b0000010100;
    pxcRom[7635] <= 10'b0000001010;
    pxcRom[7636] <= 10'b0000000101;
    pxcRom[7637] <= 10'b0000000010;
    pxcRom[7638] <= 10'b0000000001;
    pxcRom[7639] <= 10'b0000000000;
    pxcRom[7640] <= 10'b0000000000;
    pxcRom[7641] <= 10'b0000000000;
    pxcRom[7642] <= 10'b0000000000;
    pxcRom[7643] <= 10'b0000000000;
    pxcRom[7644] <= 10'b0000000000;
    pxcRom[7645] <= 10'b0000000000;
    pxcRom[7646] <= 10'b0000000000;
    pxcRom[7647] <= 10'b0000000000;
    pxcRom[7648] <= 10'b0000000000;
    pxcRom[7649] <= 10'b0000000000;
    pxcRom[7650] <= 10'b0000000000;
    pxcRom[7651] <= 10'b0000000000;
    pxcRom[7652] <= 10'b0000000001;
    pxcRom[7653] <= 10'b0000000011;
    pxcRom[7654] <= 10'b0000000111;
    pxcRom[7655] <= 10'b0000001110;
    pxcRom[7656] <= 10'b0000011001;
    pxcRom[7657] <= 10'b0000101000;
    pxcRom[7658] <= 10'b0000110001;
    pxcRom[7659] <= 10'b0000110010;
    pxcRom[7660] <= 10'b0000101000;
    pxcRom[7661] <= 10'b0000011101;
    pxcRom[7662] <= 10'b0000010010;
    pxcRom[7663] <= 10'b0000001010;
    pxcRom[7664] <= 10'b0000000101;
    pxcRom[7665] <= 10'b0000000010;
    pxcRom[7666] <= 10'b0000000001;
    pxcRom[7667] <= 10'b0000000000;
    pxcRom[7668] <= 10'b0000000000;
    pxcRom[7669] <= 10'b0000000000;
    pxcRom[7670] <= 10'b0000000000;
    pxcRom[7671] <= 10'b0000000000;
    pxcRom[7672] <= 10'b0000000000;
    pxcRom[7673] <= 10'b0000000000;
    pxcRom[7674] <= 10'b0000000000;
    pxcRom[7675] <= 10'b0000000000;
    pxcRom[7676] <= 10'b0000000000;
    pxcRom[7677] <= 10'b0000000000;
    pxcRom[7678] <= 10'b0000000000;
    pxcRom[7679] <= 10'b0000000001;
    pxcRom[7680] <= 10'b0000000010;
    pxcRom[7681] <= 10'b0000000101;
    pxcRom[7682] <= 10'b0000001011;
    pxcRom[7683] <= 10'b0000010011;
    pxcRom[7684] <= 10'b0000011111;
    pxcRom[7685] <= 10'b0000101001;
    pxcRom[7686] <= 10'b0000101100;
    pxcRom[7687] <= 10'b0000101001;
    pxcRom[7688] <= 10'b0000100001;
    pxcRom[7689] <= 10'b0000011010;
    pxcRom[7690] <= 10'b0000010001;
    pxcRom[7691] <= 10'b0000001010;
    pxcRom[7692] <= 10'b0000000101;
    pxcRom[7693] <= 10'b0000000011;
    pxcRom[7694] <= 10'b0000000001;
    pxcRom[7695] <= 10'b0000000000;
    pxcRom[7696] <= 10'b0000000000;
    pxcRom[7697] <= 10'b0000000000;
    pxcRom[7698] <= 10'b0000000000;
    pxcRom[7699] <= 10'b0000000000;
    pxcRom[7700] <= 10'b0000000000;
    pxcRom[7701] <= 10'b0000000000;
    pxcRom[7702] <= 10'b0000000000;
    pxcRom[7703] <= 10'b0000000000;
    pxcRom[7704] <= 10'b0000000000;
    pxcRom[7705] <= 10'b0000000000;
    pxcRom[7706] <= 10'b0000000000;
    pxcRom[7707] <= 10'b0000000001;
    pxcRom[7708] <= 10'b0000000100;
    pxcRom[7709] <= 10'b0000001000;
    pxcRom[7710] <= 10'b0000001111;
    pxcRom[7711] <= 10'b0000011000;
    pxcRom[7712] <= 10'b0000100001;
    pxcRom[7713] <= 10'b0000100110;
    pxcRom[7714] <= 10'b0000100110;
    pxcRom[7715] <= 10'b0000100010;
    pxcRom[7716] <= 10'b0000011101;
    pxcRom[7717] <= 10'b0000011000;
    pxcRom[7718] <= 10'b0000010000;
    pxcRom[7719] <= 10'b0000001010;
    pxcRom[7720] <= 10'b0000000110;
    pxcRom[7721] <= 10'b0000000011;
    pxcRom[7722] <= 10'b0000000001;
    pxcRom[7723] <= 10'b0000000000;
    pxcRom[7724] <= 10'b0000000000;
    pxcRom[7725] <= 10'b0000000000;
    pxcRom[7726] <= 10'b0000000000;
    pxcRom[7727] <= 10'b0000000000;
    pxcRom[7728] <= 10'b0000000000;
    pxcRom[7729] <= 10'b0000000000;
    pxcRom[7730] <= 10'b0000000000;
    pxcRom[7731] <= 10'b0000000000;
    pxcRom[7732] <= 10'b0000000000;
    pxcRom[7733] <= 10'b0000000000;
    pxcRom[7734] <= 10'b0000000001;
    pxcRom[7735] <= 10'b0000000010;
    pxcRom[7736] <= 10'b0000000101;
    pxcRom[7737] <= 10'b0000001010;
    pxcRom[7738] <= 10'b0000010001;
    pxcRom[7739] <= 10'b0000011000;
    pxcRom[7740] <= 10'b0000011111;
    pxcRom[7741] <= 10'b0000100000;
    pxcRom[7742] <= 10'b0000011111;
    pxcRom[7743] <= 10'b0000011100;
    pxcRom[7744] <= 10'b0000011001;
    pxcRom[7745] <= 10'b0000010101;
    pxcRom[7746] <= 10'b0000001111;
    pxcRom[7747] <= 10'b0000001010;
    pxcRom[7748] <= 10'b0000000110;
    pxcRom[7749] <= 10'b0000000011;
    pxcRom[7750] <= 10'b0000000001;
    pxcRom[7751] <= 10'b0000000000;
    pxcRom[7752] <= 10'b0000000000;
    pxcRom[7753] <= 10'b0000000000;
    pxcRom[7754] <= 10'b0000000000;
    pxcRom[7755] <= 10'b0000000000;
    pxcRom[7756] <= 10'b0000000000;
    pxcRom[7757] <= 10'b0000000000;
    pxcRom[7758] <= 10'b0000000000;
    pxcRom[7759] <= 10'b0000000000;
    pxcRom[7760] <= 10'b0000000000;
    pxcRom[7761] <= 10'b0000000000;
    pxcRom[7762] <= 10'b0000000001;
    pxcRom[7763] <= 10'b0000000010;
    pxcRom[7764] <= 10'b0000000100;
    pxcRom[7765] <= 10'b0000001000;
    pxcRom[7766] <= 10'b0000001110;
    pxcRom[7767] <= 10'b0000010011;
    pxcRom[7768] <= 10'b0000010111;
    pxcRom[7769] <= 10'b0000010111;
    pxcRom[7770] <= 10'b0000010110;
    pxcRom[7771] <= 10'b0000010100;
    pxcRom[7772] <= 10'b0000010010;
    pxcRom[7773] <= 10'b0000010000;
    pxcRom[7774] <= 10'b0000001100;
    pxcRom[7775] <= 10'b0000000111;
    pxcRom[7776] <= 10'b0000000100;
    pxcRom[7777] <= 10'b0000000010;
    pxcRom[7778] <= 10'b0000000001;
    pxcRom[7779] <= 10'b0000000000;
    pxcRom[7780] <= 10'b0000000000;
    pxcRom[7781] <= 10'b0000000000;
    pxcRom[7782] <= 10'b0000000000;
    pxcRom[7783] <= 10'b0000000000;
    pxcRom[7784] <= 10'b0000000000;
    pxcRom[7785] <= 10'b0000000000;
    pxcRom[7786] <= 10'b0000000000;
    pxcRom[7787] <= 10'b0000000000;
    pxcRom[7788] <= 10'b0000000000;
    pxcRom[7789] <= 10'b0000000000;
    pxcRom[7790] <= 10'b0000000000;
    pxcRom[7791] <= 10'b0000000000;
    pxcRom[7792] <= 10'b0000000001;
    pxcRom[7793] <= 10'b0000000010;
    pxcRom[7794] <= 10'b0000000011;
    pxcRom[7795] <= 10'b0000000101;
    pxcRom[7796] <= 10'b0000000110;
    pxcRom[7797] <= 10'b0000000110;
    pxcRom[7798] <= 10'b0000000110;
    pxcRom[7799] <= 10'b0000000101;
    pxcRom[7800] <= 10'b0000000100;
    pxcRom[7801] <= 10'b0000000100;
    pxcRom[7802] <= 10'b0000000011;
    pxcRom[7803] <= 10'b0000000010;
    pxcRom[7804] <= 10'b0000000001;
    pxcRom[7805] <= 10'b0000000000;
    pxcRom[7806] <= 10'b0000000000;
    pxcRom[7807] <= 10'b0000000000;
    pxcRom[7808] <= 10'b0000000000;
    pxcRom[7809] <= 10'b0000000000;
    pxcRom[7810] <= 10'b0000000000;
    pxcRom[7811] <= 10'b0000000000;
    pxcRom[7812] <= 10'b0000000000;
    pxcRom[7813] <= 10'b0000000000;
    pxcRom[7814] <= 10'b0000000000;
    pxcRom[7815] <= 10'b0000000000;
    pxcRom[7816] <= 10'b0000000000;
    pxcRom[7817] <= 10'b0000000000;
    pxcRom[7818] <= 10'b0000000000;
    pxcRom[7819] <= 10'b0000000000;
    pxcRom[7820] <= 10'b0000000000;
    pxcRom[7821] <= 10'b0000000000;
    pxcRom[7822] <= 10'b0000000000;
    pxcRom[7823] <= 10'b0000000000;
    pxcRom[7824] <= 10'b0000000000;
    pxcRom[7825] <= 10'b0000000000;
    pxcRom[7826] <= 10'b0000000000;
    pxcRom[7827] <= 10'b0000000000;
    pxcRom[7828] <= 10'b0000000000;
    pxcRom[7829] <= 10'b0000000000;
    pxcRom[7830] <= 10'b0000000000;
    pxcRom[7831] <= 10'b0000000000;
    pxcRom[7832] <= 10'b0000000000;
    pxcRom[7833] <= 10'b0000000000;
    pxcRom[7834] <= 10'b0000000000;
    pxcRom[7835] <= 10'b0000000000;
    pxcRom[7836] <= 10'b0000000000;
    pxcRom[7837] <= 10'b0000000000;
    pxcRom[7838] <= 10'b0000000000;
    pxcRom[7839] <= 10'b0000000000;
    pxcRom[7840] <= 10'b1000101011;
    pxcRom[7841] <= 10'b1000101011;
    pxcRom[7842] <= 10'b1000101011;
    pxcRom[7843] <= 10'b1000101011;
    pxcRom[7844] <= 10'b1000101011;
    pxcRom[7845] <= 10'b1000101011;
    pxcRom[7846] <= 10'b1000101011;
    pxcRom[7847] <= 10'b1000101011;
    pxcRom[7848] <= 10'b1000101011;
    pxcRom[7849] <= 10'b1000101011;
    pxcRom[7850] <= 10'b1000101011;
    pxcRom[7851] <= 10'b1000101011;
    pxcRom[7852] <= 10'b1000101011;
    pxcRom[7853] <= 10'b1000101011;
    pxcRom[7854] <= 10'b1000101011;
    pxcRom[7855] <= 10'b1000101011;
    pxcRom[7856] <= 10'b1000101011;
    pxcRom[7857] <= 10'b1000101011;
    pxcRom[7858] <= 10'b1000101011;
    pxcRom[7859] <= 10'b1000101011;
    pxcRom[7860] <= 10'b1000101011;
    pxcRom[7861] <= 10'b1000101011;
    pxcRom[7862] <= 10'b1000101011;
    pxcRom[7863] <= 10'b1000101011;
    pxcRom[7864] <= 10'b1000101011;
    pxcRom[7865] <= 10'b1000101011;
    pxcRom[7866] <= 10'b1000101011;
    pxcRom[7867] <= 10'b1000101011;
    pxcRom[7868] <= 10'b1000101011;
    pxcRom[7869] <= 10'b1000101011;
    pxcRom[7870] <= 10'b1000101011;
    pxcRom[7871] <= 10'b1000101011;
    pxcRom[7872] <= 10'b1000101011;
    pxcRom[7873] <= 10'b1000101011;
    pxcRom[7874] <= 10'b1000101011;
    pxcRom[7875] <= 10'b1000101011;
    pxcRom[7876] <= 10'b1000101011;
    pxcRom[7877] <= 10'b1000101011;
    pxcRom[7878] <= 10'b1000101011;
    pxcRom[7879] <= 10'b0111111111;
    pxcRom[7880] <= 10'b0111111111;
    pxcRom[7881] <= 10'b0111111111;
    pxcRom[7882] <= 10'b1000101011;
    pxcRom[7883] <= 10'b0111111111;
    pxcRom[7884] <= 10'b0111111111;
    pxcRom[7885] <= 10'b0111111111;
    pxcRom[7886] <= 10'b1000101011;
    pxcRom[7887] <= 10'b1000101011;
    pxcRom[7888] <= 10'b1000101011;
    pxcRom[7889] <= 10'b1000101011;
    pxcRom[7890] <= 10'b1000101011;
    pxcRom[7891] <= 10'b1000101011;
    pxcRom[7892] <= 10'b1000101011;
    pxcRom[7893] <= 10'b1000101011;
    pxcRom[7894] <= 10'b1000101011;
    pxcRom[7895] <= 10'b1000101011;
    pxcRom[7896] <= 10'b1000101011;
    pxcRom[7897] <= 10'b1000101011;
    pxcRom[7898] <= 10'b1000101011;
    pxcRom[7899] <= 10'b1000101011;
    pxcRom[7900] <= 10'b1000101011;
    pxcRom[7901] <= 10'b1000101011;
    pxcRom[7902] <= 10'b0111111111;
    pxcRom[7903] <= 10'b0111111111;
    pxcRom[7904] <= 10'b0111111111;
    pxcRom[7905] <= 10'b1000101011;
    pxcRom[7906] <= 10'b1000101011;
    pxcRom[7907] <= 10'b0111111111;
    pxcRom[7908] <= 10'b0111100101;
    pxcRom[7909] <= 10'b0111010011;
    pxcRom[7910] <= 10'b0111100101;
    pxcRom[7911] <= 10'b0111111111;
    pxcRom[7912] <= 10'b0111100101;
    pxcRom[7913] <= 10'b1000101011;
    pxcRom[7914] <= 10'b0111111111;
    pxcRom[7915] <= 10'b0111111111;
    pxcRom[7916] <= 10'b1000101011;
    pxcRom[7917] <= 10'b1000101011;
    pxcRom[7918] <= 10'b1000101011;
    pxcRom[7919] <= 10'b1000101011;
    pxcRom[7920] <= 10'b1000101011;
    pxcRom[7921] <= 10'b1000101011;
    pxcRom[7922] <= 10'b1000101011;
    pxcRom[7923] <= 10'b1000101011;
    pxcRom[7924] <= 10'b1000101011;
    pxcRom[7925] <= 10'b1000101011;
    pxcRom[7926] <= 10'b1000101011;
    pxcRom[7927] <= 10'b0111111111;
    pxcRom[7928] <= 10'b0111111111;
    pxcRom[7929] <= 10'b0111100101;
    pxcRom[7930] <= 10'b0111100101;
    pxcRom[7931] <= 10'b0111010011;
    pxcRom[7932] <= 10'b0111000100;
    pxcRom[7933] <= 10'b0110010010;
    pxcRom[7934] <= 10'b0101100110;
    pxcRom[7935] <= 10'b0100110001;
    pxcRom[7936] <= 10'b0100010101;
    pxcRom[7937] <= 10'b0100000000;
    pxcRom[7938] <= 10'b0011101110;
    pxcRom[7939] <= 10'b0011100111;
    pxcRom[7940] <= 10'b0011100101;
    pxcRom[7941] <= 10'b0011110010;
    pxcRom[7942] <= 10'b0011111110;
    pxcRom[7943] <= 10'b0100010011;
    pxcRom[7944] <= 10'b0100101100;
    pxcRom[7945] <= 10'b0101001100;
    pxcRom[7946] <= 10'b0110000011;
    pxcRom[7947] <= 10'b0110111001;
    pxcRom[7948] <= 10'b0111111111;
    pxcRom[7949] <= 10'b0111111111;
    pxcRom[7950] <= 10'b1000101011;
    pxcRom[7951] <= 10'b1000101011;
    pxcRom[7952] <= 10'b1000101011;
    pxcRom[7953] <= 10'b1000101011;
    pxcRom[7954] <= 10'b1000101011;
    pxcRom[7955] <= 10'b0111100101;
    pxcRom[7956] <= 10'b0111111111;
    pxcRom[7957] <= 10'b0111000100;
    pxcRom[7958] <= 10'b0110010010;
    pxcRom[7959] <= 10'b0101011001;
    pxcRom[7960] <= 10'b0100100011;
    pxcRom[7961] <= 10'b0011101111;
    pxcRom[7962] <= 10'b0011000001;
    pxcRom[7963] <= 10'b0010011001;
    pxcRom[7964] <= 10'b0001110101;
    pxcRom[7965] <= 10'b0001011100;
    pxcRom[7966] <= 10'b0001001011;
    pxcRom[7967] <= 10'b0001000001;
    pxcRom[7968] <= 10'b0000111111;
    pxcRom[7969] <= 10'b0001000011;
    pxcRom[7970] <= 10'b0001001111;
    pxcRom[7971] <= 10'b0001100001;
    pxcRom[7972] <= 10'b0010000001;
    pxcRom[7973] <= 10'b0010101000;
    pxcRom[7974] <= 10'b0011011010;
    pxcRom[7975] <= 10'b0100101011;
    pxcRom[7976] <= 10'b0110010010;
    pxcRom[7977] <= 10'b0111111111;
    pxcRom[7978] <= 10'b1000101011;
    pxcRom[7979] <= 10'b1000101011;
    pxcRom[7980] <= 10'b1000101011;
    pxcRom[7981] <= 10'b1000101011;
    pxcRom[7982] <= 10'b1000101011;
    pxcRom[7983] <= 10'b0111010011;
    pxcRom[7984] <= 10'b0111010011;
    pxcRom[7985] <= 10'b0110010010;
    pxcRom[7986] <= 10'b0101010010;
    pxcRom[7987] <= 10'b0100010101;
    pxcRom[7988] <= 10'b0011010111;
    pxcRom[7989] <= 10'b0010100101;
    pxcRom[7990] <= 10'b0001111011;
    pxcRom[7991] <= 10'b0001011000;
    pxcRom[7992] <= 10'b0000111100;
    pxcRom[7993] <= 10'b0000101001;
    pxcRom[7994] <= 10'b0000011101;
    pxcRom[7995] <= 10'b0000010110;
    pxcRom[7996] <= 10'b0000010100;
    pxcRom[7997] <= 10'b0000010111;
    pxcRom[7998] <= 10'b0000100000;
    pxcRom[7999] <= 10'b0000101111;
    pxcRom[8000] <= 10'b0001000111;
    pxcRom[8001] <= 10'b0001101001;
    pxcRom[8002] <= 10'b0010011101;
    pxcRom[8003] <= 10'b0011011111;
    pxcRom[8004] <= 10'b0101100000;
    pxcRom[8005] <= 10'b0111111111;
    pxcRom[8006] <= 10'b1000101011;
    pxcRom[8007] <= 10'b1000101011;
    pxcRom[8008] <= 10'b1000101011;
    pxcRom[8009] <= 10'b1000101011;
    pxcRom[8010] <= 10'b1000101011;
    pxcRom[8011] <= 10'b1000101011;
    pxcRom[8012] <= 10'b0110011000;
    pxcRom[8013] <= 10'b0101010100;
    pxcRom[8014] <= 10'b0100011100;
    pxcRom[8015] <= 10'b0011011100;
    pxcRom[8016] <= 10'b0010100101;
    pxcRom[8017] <= 10'b0001110110;
    pxcRom[8018] <= 10'b0001010001;
    pxcRom[8019] <= 10'b0000110100;
    pxcRom[8020] <= 10'b0000100010;
    pxcRom[8021] <= 10'b0000010101;
    pxcRom[8022] <= 10'b0000001110;
    pxcRom[8023] <= 10'b0000001010;
    pxcRom[8024] <= 10'b0000001001;
    pxcRom[8025] <= 10'b0000001010;
    pxcRom[8026] <= 10'b0000001110;
    pxcRom[8027] <= 10'b0000011000;
    pxcRom[8028] <= 10'b0000101010;
    pxcRom[8029] <= 10'b0001000011;
    pxcRom[8030] <= 10'b0001101100;
    pxcRom[8031] <= 10'b0010101000;
    pxcRom[8032] <= 10'b0100100001;
    pxcRom[8033] <= 10'b0111000100;
    pxcRom[8034] <= 10'b0111111111;
    pxcRom[8035] <= 10'b0111111111;
    pxcRom[8036] <= 10'b1000101011;
    pxcRom[8037] <= 10'b1000101011;
    pxcRom[8038] <= 10'b1000101011;
    pxcRom[8039] <= 10'b0111111111;
    pxcRom[8040] <= 10'b0110011000;
    pxcRom[8041] <= 10'b0100110010;
    pxcRom[8042] <= 10'b0011110001;
    pxcRom[8043] <= 10'b0010101100;
    pxcRom[8044] <= 10'b0001110111;
    pxcRom[8045] <= 10'b0001010001;
    pxcRom[8046] <= 10'b0000110100;
    pxcRom[8047] <= 10'b0000100000;
    pxcRom[8048] <= 10'b0000010100;
    pxcRom[8049] <= 10'b0000001101;
    pxcRom[8050] <= 10'b0000001011;
    pxcRom[8051] <= 10'b0000001010;
    pxcRom[8052] <= 10'b0000001001;
    pxcRom[8053] <= 10'b0000001000;
    pxcRom[8054] <= 10'b0000001001;
    pxcRom[8055] <= 10'b0000001110;
    pxcRom[8056] <= 10'b0000011001;
    pxcRom[8057] <= 10'b0000101101;
    pxcRom[8058] <= 10'b0001001100;
    pxcRom[8059] <= 10'b0010000000;
    pxcRom[8060] <= 10'b0011101000;
    pxcRom[8061] <= 10'b0110100110;
    pxcRom[8062] <= 10'b1000101011;
    pxcRom[8063] <= 10'b0111111111;
    pxcRom[8064] <= 10'b0111111111;
    pxcRom[8065] <= 10'b1000101011;
    pxcRom[8066] <= 10'b0111100101;
    pxcRom[8067] <= 10'b0111010011;
    pxcRom[8068] <= 10'b0110000011;
    pxcRom[8069] <= 10'b0100011010;
    pxcRom[8070] <= 10'b0011000011;
    pxcRom[8071] <= 10'b0010000100;
    pxcRom[8072] <= 10'b0001010111;
    pxcRom[8073] <= 10'b0000111000;
    pxcRom[8074] <= 10'b0000100001;
    pxcRom[8075] <= 10'b0000010101;
    pxcRom[8076] <= 10'b0000001111;
    pxcRom[8077] <= 10'b0000001110;
    pxcRom[8078] <= 10'b0000010000;
    pxcRom[8079] <= 10'b0000010011;
    pxcRom[8080] <= 10'b0000010100;
    pxcRom[8081] <= 10'b0000010001;
    pxcRom[8082] <= 10'b0000001110;
    pxcRom[8083] <= 10'b0000001100;
    pxcRom[8084] <= 10'b0000010001;
    pxcRom[8085] <= 10'b0000011110;
    pxcRom[8086] <= 10'b0000111000;
    pxcRom[8087] <= 10'b0001100011;
    pxcRom[8088] <= 10'b0010111101;
    pxcRom[8089] <= 10'b0110100110;
    pxcRom[8090] <= 10'b1000101011;
    pxcRom[8091] <= 10'b1000101011;
    pxcRom[8092] <= 10'b1000101011;
    pxcRom[8093] <= 10'b1000101011;
    pxcRom[8094] <= 10'b1000101011;
    pxcRom[8095] <= 10'b0111111111;
    pxcRom[8096] <= 10'b0101101111;
    pxcRom[8097] <= 10'b0011101010;
    pxcRom[8098] <= 10'b0010011100;
    pxcRom[8099] <= 10'b0001100011;
    pxcRom[8100] <= 10'b0000111111;
    pxcRom[8101] <= 10'b0000100101;
    pxcRom[8102] <= 10'b0000010110;
    pxcRom[8103] <= 10'b0000010000;
    pxcRom[8104] <= 10'b0000010000;
    pxcRom[8105] <= 10'b0000010101;
    pxcRom[8106] <= 10'b0000011110;
    pxcRom[8107] <= 10'b0000100101;
    pxcRom[8108] <= 10'b0000101000;
    pxcRom[8109] <= 10'b0000100110;
    pxcRom[8110] <= 10'b0000011100;
    pxcRom[8111] <= 10'b0000010010;
    pxcRom[8112] <= 10'b0000001111;
    pxcRom[8113] <= 10'b0000010110;
    pxcRom[8114] <= 10'b0000101010;
    pxcRom[8115] <= 10'b0001001110;
    pxcRom[8116] <= 10'b0010100011;
    pxcRom[8117] <= 10'b0110011000;
    pxcRom[8118] <= 10'b1000101011;
    pxcRom[8119] <= 10'b1000101011;
    pxcRom[8120] <= 10'b1000101011;
    pxcRom[8121] <= 10'b1000101011;
    pxcRom[8122] <= 10'b0111111111;
    pxcRom[8123] <= 10'b0111100101;
    pxcRom[8124] <= 10'b0101001000;
    pxcRom[8125] <= 10'b0010111111;
    pxcRom[8126] <= 10'b0001111001;
    pxcRom[8127] <= 10'b0001001010;
    pxcRom[8128] <= 10'b0000101100;
    pxcRom[8129] <= 10'b0000011001;
    pxcRom[8130] <= 10'b0000010000;
    pxcRom[8131] <= 10'b0000010000;
    pxcRom[8132] <= 10'b0000011000;
    pxcRom[8133] <= 10'b0000100100;
    pxcRom[8134] <= 10'b0000110010;
    pxcRom[8135] <= 10'b0001000010;
    pxcRom[8136] <= 10'b0001001010;
    pxcRom[8137] <= 10'b0001000100;
    pxcRom[8138] <= 10'b0000101111;
    pxcRom[8139] <= 10'b0000011011;
    pxcRom[8140] <= 10'b0000010001;
    pxcRom[8141] <= 10'b0000010010;
    pxcRom[8142] <= 10'b0000100001;
    pxcRom[8143] <= 10'b0000111111;
    pxcRom[8144] <= 10'b0010001100;
    pxcRom[8145] <= 10'b0110000011;
    pxcRom[8146] <= 10'b1000101011;
    pxcRom[8147] <= 10'b1000101011;
    pxcRom[8148] <= 10'b1000101011;
    pxcRom[8149] <= 10'b0111111111;
    pxcRom[8150] <= 10'b1000101011;
    pxcRom[8151] <= 10'b0111111111;
    pxcRom[8152] <= 10'b0100100011;
    pxcRom[8153] <= 10'b0010011010;
    pxcRom[8154] <= 10'b0001011101;
    pxcRom[8155] <= 10'b0000110111;
    pxcRom[8156] <= 10'b0000011111;
    pxcRom[8157] <= 10'b0000010010;
    pxcRom[8158] <= 10'b0000001111;
    pxcRom[8159] <= 10'b0000010110;
    pxcRom[8160] <= 10'b0000100101;
    pxcRom[8161] <= 10'b0000111001;
    pxcRom[8162] <= 10'b0001010001;
    pxcRom[8163] <= 10'b0001101001;
    pxcRom[8164] <= 10'b0001110011;
    pxcRom[8165] <= 10'b0001100011;
    pxcRom[8166] <= 10'b0001000011;
    pxcRom[8167] <= 10'b0000100110;
    pxcRom[8168] <= 10'b0000010100;
    pxcRom[8169] <= 10'b0000010000;
    pxcRom[8170] <= 10'b0000011011;
    pxcRom[8171] <= 10'b0000110110;
    pxcRom[8172] <= 10'b0001111010;
    pxcRom[8173] <= 10'b0101011011;
    pxcRom[8174] <= 10'b0111111111;
    pxcRom[8175] <= 10'b1000101011;
    pxcRom[8176] <= 10'b1000101011;
    pxcRom[8177] <= 10'b1000101011;
    pxcRom[8178] <= 10'b0111111111;
    pxcRom[8179] <= 10'b0111111111;
    pxcRom[8180] <= 10'b0011110110;
    pxcRom[8181] <= 10'b0001111100;
    pxcRom[8182] <= 10'b0001001000;
    pxcRom[8183] <= 10'b0000100111;
    pxcRom[8184] <= 10'b0000010101;
    pxcRom[8185] <= 10'b0000001111;
    pxcRom[8186] <= 10'b0000010011;
    pxcRom[8187] <= 10'b0000100010;
    pxcRom[8188] <= 10'b0000111001;
    pxcRom[8189] <= 10'b0001011000;
    pxcRom[8190] <= 10'b0001111101;
    pxcRom[8191] <= 10'b0010011001;
    pxcRom[8192] <= 10'b0010011010;
    pxcRom[8193] <= 10'b0001111011;
    pxcRom[8194] <= 10'b0001010000;
    pxcRom[8195] <= 10'b0000101101;
    pxcRom[8196] <= 10'b0000010111;
    pxcRom[8197] <= 10'b0000010001;
    pxcRom[8198] <= 10'b0000011001;
    pxcRom[8199] <= 10'b0000110010;
    pxcRom[8200] <= 10'b0001101111;
    pxcRom[8201] <= 10'b0101000100;
    pxcRom[8202] <= 10'b0111111111;
    pxcRom[8203] <= 10'b1000101011;
    pxcRom[8204] <= 10'b1000101011;
    pxcRom[8205] <= 10'b0111111111;
    pxcRom[8206] <= 10'b0111100101;
    pxcRom[8207] <= 10'b0111010011;
    pxcRom[8208] <= 10'b0011010110;
    pxcRom[8209] <= 10'b0001100011;
    pxcRom[8210] <= 10'b0000110110;
    pxcRom[8211] <= 10'b0000011100;
    pxcRom[8212] <= 10'b0000010000;
    pxcRom[8213] <= 10'b0000010000;
    pxcRom[8214] <= 10'b0000011011;
    pxcRom[8215] <= 10'b0000110010;
    pxcRom[8216] <= 10'b0001010110;
    pxcRom[8217] <= 10'b0010000011;
    pxcRom[8218] <= 10'b0010110000;
    pxcRom[8219] <= 10'b0011000111;
    pxcRom[8220] <= 10'b0010111101;
    pxcRom[8221] <= 10'b0010000101;
    pxcRom[8222] <= 10'b0001010011;
    pxcRom[8223] <= 10'b0000101111;
    pxcRom[8224] <= 10'b0000011000;
    pxcRom[8225] <= 10'b0000010001;
    pxcRom[8226] <= 10'b0000011010;
    pxcRom[8227] <= 10'b0000110010;
    pxcRom[8228] <= 10'b0001101101;
    pxcRom[8229] <= 10'b0100111011;
    pxcRom[8230] <= 10'b1000101011;
    pxcRom[8231] <= 10'b1000101011;
    pxcRom[8232] <= 10'b1000101011;
    pxcRom[8233] <= 10'b1000101011;
    pxcRom[8234] <= 10'b1000101011;
    pxcRom[8235] <= 10'b0111100101;
    pxcRom[8236] <= 10'b0010110110;
    pxcRom[8237] <= 10'b0001010000;
    pxcRom[8238] <= 10'b0000101010;
    pxcRom[8239] <= 10'b0000010101;
    pxcRom[8240] <= 10'b0000001111;
    pxcRom[8241] <= 10'b0000010100;
    pxcRom[8242] <= 10'b0000100111;
    pxcRom[8243] <= 10'b0001001000;
    pxcRom[8244] <= 10'b0001111010;
    pxcRom[8245] <= 10'b0010110001;
    pxcRom[8246] <= 10'b0011011011;
    pxcRom[8247] <= 10'b0011101001;
    pxcRom[8248] <= 10'b0010111110;
    pxcRom[8249] <= 10'b0001111110;
    pxcRom[8250] <= 10'b0001001110;
    pxcRom[8251] <= 10'b0000101011;
    pxcRom[8252] <= 10'b0000010111;
    pxcRom[8253] <= 10'b0000010010;
    pxcRom[8254] <= 10'b0000011100;
    pxcRom[8255] <= 10'b0000110110;
    pxcRom[8256] <= 10'b0001101111;
    pxcRom[8257] <= 10'b0100110001;
    pxcRom[8258] <= 10'b1000101011;
    pxcRom[8259] <= 10'b1000101011;
    pxcRom[8260] <= 10'b1000101011;
    pxcRom[8261] <= 10'b1000101011;
    pxcRom[8262] <= 10'b1000101011;
    pxcRom[8263] <= 10'b0111010011;
    pxcRom[8264] <= 10'b0010011011;
    pxcRom[8265] <= 10'b0001000001;
    pxcRom[8266] <= 10'b0000100001;
    pxcRom[8267] <= 10'b0000010001;
    pxcRom[8268] <= 10'b0000001111;
    pxcRom[8269] <= 10'b0000011010;
    pxcRom[8270] <= 10'b0000110011;
    pxcRom[8271] <= 10'b0001100010;
    pxcRom[8272] <= 10'b0010011101;
    pxcRom[8273] <= 10'b0011011000;
    pxcRom[8274] <= 10'b0011111001;
    pxcRom[8275] <= 10'b0011011100;
    pxcRom[8276] <= 10'b0010100101;
    pxcRom[8277] <= 10'b0001101001;
    pxcRom[8278] <= 10'b0001000000;
    pxcRom[8279] <= 10'b0000100100;
    pxcRom[8280] <= 10'b0000010101;
    pxcRom[8281] <= 10'b0000010100;
    pxcRom[8282] <= 10'b0000100000;
    pxcRom[8283] <= 10'b0000111101;
    pxcRom[8284] <= 10'b0001110111;
    pxcRom[8285] <= 10'b0100101101;
    pxcRom[8286] <= 10'b1000101011;
    pxcRom[8287] <= 10'b1000101011;
    pxcRom[8288] <= 10'b1000101011;
    pxcRom[8289] <= 10'b1000101011;
    pxcRom[8290] <= 10'b1000101011;
    pxcRom[8291] <= 10'b0110100110;
    pxcRom[8292] <= 10'b0010001010;
    pxcRom[8293] <= 10'b0000110111;
    pxcRom[8294] <= 10'b0000011100;
    pxcRom[8295] <= 10'b0000001111;
    pxcRom[8296] <= 10'b0000010000;
    pxcRom[8297] <= 10'b0000100001;
    pxcRom[8298] <= 10'b0001000001;
    pxcRom[8299] <= 10'b0001110111;
    pxcRom[8300] <= 10'b0010110101;
    pxcRom[8301] <= 10'b0011101010;
    pxcRom[8302] <= 10'b0011100100;
    pxcRom[8303] <= 10'b0010110000;
    pxcRom[8304] <= 10'b0001111011;
    pxcRom[8305] <= 10'b0001001111;
    pxcRom[8306] <= 10'b0000101111;
    pxcRom[8307] <= 10'b0000011011;
    pxcRom[8308] <= 10'b0000010011;
    pxcRom[8309] <= 10'b0000011000;
    pxcRom[8310] <= 10'b0000101000;
    pxcRom[8311] <= 10'b0001000111;
    pxcRom[8312] <= 10'b0010000110;
    pxcRom[8313] <= 10'b0101000001;
    pxcRom[8314] <= 10'b1000101011;
    pxcRom[8315] <= 10'b1000101011;
    pxcRom[8316] <= 10'b1000101011;
    pxcRom[8317] <= 10'b1000101011;
    pxcRom[8318] <= 10'b1000101011;
    pxcRom[8319] <= 10'b0110011111;
    pxcRom[8320] <= 10'b0001111110;
    pxcRom[8321] <= 10'b0000110011;
    pxcRom[8322] <= 10'b0000011010;
    pxcRom[8323] <= 10'b0000001110;
    pxcRom[8324] <= 10'b0000010001;
    pxcRom[8325] <= 10'b0000100101;
    pxcRom[8326] <= 10'b0001001000;
    pxcRom[8327] <= 10'b0001111101;
    pxcRom[8328] <= 10'b0010101110;
    pxcRom[8329] <= 10'b0010111100;
    pxcRom[8330] <= 10'b0010100011;
    pxcRom[8331] <= 10'b0001111010;
    pxcRom[8332] <= 10'b0001010100;
    pxcRom[8333] <= 10'b0000110011;
    pxcRom[8334] <= 10'b0000100000;
    pxcRom[8335] <= 10'b0000010100;
    pxcRom[8336] <= 10'b0000010011;
    pxcRom[8337] <= 10'b0000011110;
    pxcRom[8338] <= 10'b0000110110;
    pxcRom[8339] <= 10'b0001011011;
    pxcRom[8340] <= 10'b0010011100;
    pxcRom[8341] <= 10'b0101100110;
    pxcRom[8342] <= 10'b1000101011;
    pxcRom[8343] <= 10'b0111111111;
    pxcRom[8344] <= 10'b1000101011;
    pxcRom[8345] <= 10'b1000101011;
    pxcRom[8346] <= 10'b1000101011;
    pxcRom[8347] <= 10'b0110001100;
    pxcRom[8348] <= 10'b0001111001;
    pxcRom[8349] <= 10'b0000110100;
    pxcRom[8350] <= 10'b0000011010;
    pxcRom[8351] <= 10'b0000001110;
    pxcRom[8352] <= 10'b0000010001;
    pxcRom[8353] <= 10'b0000100010;
    pxcRom[8354] <= 10'b0001000000;
    pxcRom[8355] <= 10'b0001100101;
    pxcRom[8356] <= 10'b0001111110;
    pxcRom[8357] <= 10'b0001111011;
    pxcRom[8358] <= 10'b0001100100;
    pxcRom[8359] <= 10'b0001001001;
    pxcRom[8360] <= 10'b0000110001;
    pxcRom[8361] <= 10'b0000100000;
    pxcRom[8362] <= 10'b0000010101;
    pxcRom[8363] <= 10'b0000010010;
    pxcRom[8364] <= 10'b0000011001;
    pxcRom[8365] <= 10'b0000101011;
    pxcRom[8366] <= 10'b0001000111;
    pxcRom[8367] <= 10'b0001110101;
    pxcRom[8368] <= 10'b0011000010;
    pxcRom[8369] <= 10'b0110000111;
    pxcRom[8370] <= 10'b1000101011;
    pxcRom[8371] <= 10'b1000101011;
    pxcRom[8372] <= 10'b1000101011;
    pxcRom[8373] <= 10'b0111111111;
    pxcRom[8374] <= 10'b0111111111;
    pxcRom[8375] <= 10'b0101110010;
    pxcRom[8376] <= 10'b0001111100;
    pxcRom[8377] <= 10'b0000111000;
    pxcRom[8378] <= 10'b0000011101;
    pxcRom[8379] <= 10'b0000001111;
    pxcRom[8380] <= 10'b0000001110;
    pxcRom[8381] <= 10'b0000011000;
    pxcRom[8382] <= 10'b0000101010;
    pxcRom[8383] <= 10'b0000111110;
    pxcRom[8384] <= 10'b0001000111;
    pxcRom[8385] <= 10'b0001000100;
    pxcRom[8386] <= 10'b0000110111;
    pxcRom[8387] <= 10'b0000101000;
    pxcRom[8388] <= 10'b0000011011;
    pxcRom[8389] <= 10'b0000010011;
    pxcRom[8390] <= 10'b0000010000;
    pxcRom[8391] <= 10'b0000010101;
    pxcRom[8392] <= 10'b0000100101;
    pxcRom[8393] <= 10'b0000111110;
    pxcRom[8394] <= 10'b0001100010;
    pxcRom[8395] <= 10'b0010011010;
    pxcRom[8396] <= 10'b0011110111;
    pxcRom[8397] <= 10'b0110111001;
    pxcRom[8398] <= 10'b1000101011;
    pxcRom[8399] <= 10'b1000101011;
    pxcRom[8400] <= 10'b1000101011;
    pxcRom[8401] <= 10'b0111111111;
    pxcRom[8402] <= 10'b0111111111;
    pxcRom[8403] <= 10'b0101110110;
    pxcRom[8404] <= 10'b0010001011;
    pxcRom[8405] <= 10'b0001000101;
    pxcRom[8406] <= 10'b0000100100;
    pxcRom[8407] <= 10'b0000010010;
    pxcRom[8408] <= 10'b0000001011;
    pxcRom[8409] <= 10'b0000001101;
    pxcRom[8410] <= 10'b0000010100;
    pxcRom[8411] <= 10'b0000011100;
    pxcRom[8412] <= 10'b0000011111;
    pxcRom[8413] <= 10'b0000011111;
    pxcRom[8414] <= 10'b0000011001;
    pxcRom[8415] <= 10'b0000010011;
    pxcRom[8416] <= 10'b0000001111;
    pxcRom[8417] <= 10'b0000001111;
    pxcRom[8418] <= 10'b0000010101;
    pxcRom[8419] <= 10'b0000100100;
    pxcRom[8420] <= 10'b0000111010;
    pxcRom[8421] <= 10'b0001011001;
    pxcRom[8422] <= 10'b0010001011;
    pxcRom[8423] <= 10'b0011010000;
    pxcRom[8424] <= 10'b0100111001;
    pxcRom[8425] <= 10'b0111100101;
    pxcRom[8426] <= 10'b0111111111;
    pxcRom[8427] <= 10'b1000101011;
    pxcRom[8428] <= 10'b1000101011;
    pxcRom[8429] <= 10'b1000101011;
    pxcRom[8430] <= 10'b0111111111;
    pxcRom[8431] <= 10'b0101111110;
    pxcRom[8432] <= 10'b0010100011;
    pxcRom[8433] <= 10'b0001011100;
    pxcRom[8434] <= 10'b0000110011;
    pxcRom[8435] <= 10'b0000011011;
    pxcRom[8436] <= 10'b0000001101;
    pxcRom[8437] <= 10'b0000001000;
    pxcRom[8438] <= 10'b0000000111;
    pxcRom[8439] <= 10'b0000001001;
    pxcRom[8440] <= 10'b0000001011;
    pxcRom[8441] <= 10'b0000001100;
    pxcRom[8442] <= 10'b0000001011;
    pxcRom[8443] <= 10'b0000001011;
    pxcRom[8444] <= 10'b0000001110;
    pxcRom[8445] <= 10'b0000010110;
    pxcRom[8446] <= 10'b0000100110;
    pxcRom[8447] <= 10'b0000111100;
    pxcRom[8448] <= 10'b0001011011;
    pxcRom[8449] <= 10'b0010000111;
    pxcRom[8450] <= 10'b0011000100;
    pxcRom[8451] <= 10'b0100010111;
    pxcRom[8452] <= 10'b0101111010;
    pxcRom[8453] <= 10'b0111111111;
    pxcRom[8454] <= 10'b0111010011;
    pxcRom[8455] <= 10'b0111111111;
    pxcRom[8456] <= 10'b1000101011;
    pxcRom[8457] <= 10'b1000101011;
    pxcRom[8458] <= 10'b1000101011;
    pxcRom[8459] <= 10'b0110100110;
    pxcRom[8460] <= 10'b0011011000;
    pxcRom[8461] <= 10'b0010000000;
    pxcRom[8462] <= 10'b0001001111;
    pxcRom[8463] <= 10'b0000101111;
    pxcRom[8464] <= 10'b0000011010;
    pxcRom[8465] <= 10'b0000001110;
    pxcRom[8466] <= 10'b0000001000;
    pxcRom[8467] <= 10'b0000000111;
    pxcRom[8468] <= 10'b0000000111;
    pxcRom[8469] <= 10'b0000001000;
    pxcRom[8470] <= 10'b0000001011;
    pxcRom[8471] <= 10'b0000010010;
    pxcRom[8472] <= 10'b0000011101;
    pxcRom[8473] <= 10'b0000101110;
    pxcRom[8474] <= 10'b0001000110;
    pxcRom[8475] <= 10'b0001100110;
    pxcRom[8476] <= 10'b0010010010;
    pxcRom[8477] <= 10'b0011001101;
    pxcRom[8478] <= 10'b0100010110;
    pxcRom[8479] <= 10'b0101101111;
    pxcRom[8480] <= 10'b0110101111;
    pxcRom[8481] <= 10'b0111010011;
    pxcRom[8482] <= 10'b0111111111;
    pxcRom[8483] <= 10'b0111111111;
    pxcRom[8484] <= 10'b1000101011;
    pxcRom[8485] <= 10'b1000101011;
    pxcRom[8486] <= 10'b1000101011;
    pxcRom[8487] <= 10'b0111111111;
    pxcRom[8488] <= 10'b0100110010;
    pxcRom[8489] <= 10'b0011000101;
    pxcRom[8490] <= 10'b0010000100;
    pxcRom[8491] <= 10'b0001011000;
    pxcRom[8492] <= 10'b0000111010;
    pxcRom[8493] <= 10'b0000100111;
    pxcRom[8494] <= 10'b0000011010;
    pxcRom[8495] <= 10'b0000010101;
    pxcRom[8496] <= 10'b0000010100;
    pxcRom[8497] <= 10'b0000011000;
    pxcRom[8498] <= 10'b0000100001;
    pxcRom[8499] <= 10'b0000101111;
    pxcRom[8500] <= 10'b0001000001;
    pxcRom[8501] <= 10'b0001011100;
    pxcRom[8502] <= 10'b0001111111;
    pxcRom[8503] <= 10'b0010101111;
    pxcRom[8504] <= 10'b0011101101;
    pxcRom[8505] <= 10'b0100111011;
    pxcRom[8506] <= 10'b0101110010;
    pxcRom[8507] <= 10'b0110011111;
    pxcRom[8508] <= 10'b0111000100;
    pxcRom[8509] <= 10'b0111100101;
    pxcRom[8510] <= 10'b1000101011;
    pxcRom[8511] <= 10'b1000101011;
    pxcRom[8512] <= 10'b1000101011;
    pxcRom[8513] <= 10'b1000101011;
    pxcRom[8514] <= 10'b1000101011;
    pxcRom[8515] <= 10'b1000101011;
    pxcRom[8516] <= 10'b0110100110;
    pxcRom[8517] <= 10'b0101010000;
    pxcRom[8518] <= 10'b0100000000;
    pxcRom[8519] <= 10'b0011001000;
    pxcRom[8520] <= 10'b0010100000;
    pxcRom[8521] <= 10'b0010000011;
    pxcRom[8522] <= 10'b0001110010;
    pxcRom[8523] <= 10'b0001101000;
    pxcRom[8524] <= 10'b0001100100;
    pxcRom[8525] <= 10'b0001101001;
    pxcRom[8526] <= 10'b0001110100;
    pxcRom[8527] <= 10'b0010000110;
    pxcRom[8528] <= 10'b0010100001;
    pxcRom[8529] <= 10'b0011000011;
    pxcRom[8530] <= 10'b0011110101;
    pxcRom[8531] <= 10'b0100101011;
    pxcRom[8532] <= 10'b0101101111;
    pxcRom[8533] <= 10'b0111000100;
    pxcRom[8534] <= 10'b0111000100;
    pxcRom[8535] <= 10'b0111100101;
    pxcRom[8536] <= 10'b0111100101;
    pxcRom[8537] <= 10'b0111111111;
    pxcRom[8538] <= 10'b1000101011;
    pxcRom[8539] <= 10'b1000101011;
    pxcRom[8540] <= 10'b1000101011;
    pxcRom[8541] <= 10'b1000101011;
    pxcRom[8542] <= 10'b1000101011;
    pxcRom[8543] <= 10'b1000101011;
    pxcRom[8544] <= 10'b1000101011;
    pxcRom[8545] <= 10'b1000101011;
    pxcRom[8546] <= 10'b0111111111;
    pxcRom[8547] <= 10'b0111100101;
    pxcRom[8548] <= 10'b0110100110;
    pxcRom[8549] <= 10'b0101111110;
    pxcRom[8550] <= 10'b0101110110;
    pxcRom[8551] <= 10'b0101101111;
    pxcRom[8552] <= 10'b0101110010;
    pxcRom[8553] <= 10'b0101111110;
    pxcRom[8554] <= 10'b0110000111;
    pxcRom[8555] <= 10'b0110100110;
    pxcRom[8556] <= 10'b0111000100;
    pxcRom[8557] <= 10'b0111111111;
    pxcRom[8558] <= 10'b0111111111;
    pxcRom[8559] <= 10'b1000101011;
    pxcRom[8560] <= 10'b1000101011;
    pxcRom[8561] <= 10'b1000101011;
    pxcRom[8562] <= 10'b1000101011;
    pxcRom[8563] <= 10'b1000101011;
    pxcRom[8564] <= 10'b1000101011;
    pxcRom[8565] <= 10'b1000101011;
    pxcRom[8566] <= 10'b1000101011;
    pxcRom[8567] <= 10'b1000101011;
    pxcRom[8568] <= 10'b1000101011;
    pxcRom[8569] <= 10'b1000101011;
    pxcRom[8570] <= 10'b1000101011;
    pxcRom[8571] <= 10'b1000101011;
    pxcRom[8572] <= 10'b1000101011;
    pxcRom[8573] <= 10'b1000101011;
    pxcRom[8574] <= 10'b1000101011;
    pxcRom[8575] <= 10'b1000101011;
    pxcRom[8576] <= 10'b1000101011;
    pxcRom[8577] <= 10'b1000101011;
    pxcRom[8578] <= 10'b1000101011;
    pxcRom[8579] <= 10'b1000101011;
    pxcRom[8580] <= 10'b1000101011;
    pxcRom[8581] <= 10'b1000101011;
    pxcRom[8582] <= 10'b1000101011;
    pxcRom[8583] <= 10'b1000101011;
    pxcRom[8584] <= 10'b1000101011;
    pxcRom[8585] <= 10'b1000101011;
    pxcRom[8586] <= 10'b1000101011;
    pxcRom[8587] <= 10'b1000101011;
    pxcRom[8588] <= 10'b1000101011;
    pxcRom[8589] <= 10'b1000101011;
    pxcRom[8590] <= 10'b1000101011;
    pxcRom[8591] <= 10'b1000101011;
    pxcRom[8592] <= 10'b1000101011;
    pxcRom[8593] <= 10'b1000101011;
    pxcRom[8594] <= 10'b1000101011;
    pxcRom[8595] <= 10'b1000101011;
    pxcRom[8596] <= 10'b1000101011;
    pxcRom[8597] <= 10'b1000101011;
    pxcRom[8598] <= 10'b1000101011;
    pxcRom[8599] <= 10'b1000101011;
    pxcRom[8600] <= 10'b1000101011;
    pxcRom[8601] <= 10'b1000101011;
    pxcRom[8602] <= 10'b1000101011;
    pxcRom[8603] <= 10'b1000101011;
    pxcRom[8604] <= 10'b1000101011;
    pxcRom[8605] <= 10'b1000101011;
    pxcRom[8606] <= 10'b1000101011;
    pxcRom[8607] <= 10'b1000101011;
    pxcRom[8608] <= 10'b1000101011;
    pxcRom[8609] <= 10'b1000101011;
    pxcRom[8610] <= 10'b1000101011;
    pxcRom[8611] <= 10'b1000101011;
    pxcRom[8612] <= 10'b1000101011;
    pxcRom[8613] <= 10'b1000101011;
    pxcRom[8614] <= 10'b1000101011;
    pxcRom[8615] <= 10'b1000101011;
    pxcRom[8616] <= 10'b1000101011;
    pxcRom[8617] <= 10'b1000101011;
    pxcRom[8618] <= 10'b1000101011;
    pxcRom[8619] <= 10'b1000101011;
    pxcRom[8620] <= 10'b1000101011;
    pxcRom[8621] <= 10'b1000101011;
    pxcRom[8622] <= 10'b1000101011;
    pxcRom[8623] <= 10'b1000101011;
    pxcRom[8624] <= 10'b1000110100;
    pxcRom[8625] <= 10'b1000110100;
    pxcRom[8626] <= 10'b1000110100;
    pxcRom[8627] <= 10'b1000110100;
    pxcRom[8628] <= 10'b1000110100;
    pxcRom[8629] <= 10'b1000110100;
    pxcRom[8630] <= 10'b1000110100;
    pxcRom[8631] <= 10'b1000110100;
    pxcRom[8632] <= 10'b1000110100;
    pxcRom[8633] <= 10'b1000110100;
    pxcRom[8634] <= 10'b1000110100;
    pxcRom[8635] <= 10'b1000110100;
    pxcRom[8636] <= 10'b1000110100;
    pxcRom[8637] <= 10'b1000110100;
    pxcRom[8638] <= 10'b1000110100;
    pxcRom[8639] <= 10'b1000110100;
    pxcRom[8640] <= 10'b1000110100;
    pxcRom[8641] <= 10'b1000110100;
    pxcRom[8642] <= 10'b1000110100;
    pxcRom[8643] <= 10'b1000110100;
    pxcRom[8644] <= 10'b1000110100;
    pxcRom[8645] <= 10'b1000110100;
    pxcRom[8646] <= 10'b1000110100;
    pxcRom[8647] <= 10'b1000110100;
    pxcRom[8648] <= 10'b1000110100;
    pxcRom[8649] <= 10'b1000110100;
    pxcRom[8650] <= 10'b1000110100;
    pxcRom[8651] <= 10'b1000110100;
    pxcRom[8652] <= 10'b1000110100;
    pxcRom[8653] <= 10'b1000110100;
    pxcRom[8654] <= 10'b1000110100;
    pxcRom[8655] <= 10'b1000110100;
    pxcRom[8656] <= 10'b1000110100;
    pxcRom[8657] <= 10'b1000110100;
    pxcRom[8658] <= 10'b1000110100;
    pxcRom[8659] <= 10'b1000110100;
    pxcRom[8660] <= 10'b1000110100;
    pxcRom[8661] <= 10'b1000110100;
    pxcRom[8662] <= 10'b1000110100;
    pxcRom[8663] <= 10'b1000110100;
    pxcRom[8664] <= 10'b1000110100;
    pxcRom[8665] <= 10'b1000110100;
    pxcRom[8666] <= 10'b0111101101;
    pxcRom[8667] <= 10'b0111101101;
    pxcRom[8668] <= 10'b0111101101;
    pxcRom[8669] <= 10'b1000110100;
    pxcRom[8670] <= 10'b1000110100;
    pxcRom[8671] <= 10'b1000110100;
    pxcRom[8672] <= 10'b1000110100;
    pxcRom[8673] <= 10'b1000110100;
    pxcRom[8674] <= 10'b1000110100;
    pxcRom[8675] <= 10'b1000110100;
    pxcRom[8676] <= 10'b1000110100;
    pxcRom[8677] <= 10'b1000110100;
    pxcRom[8678] <= 10'b1000110100;
    pxcRom[8679] <= 10'b1000110100;
    pxcRom[8680] <= 10'b1000110100;
    pxcRom[8681] <= 10'b1000110100;
    pxcRom[8682] <= 10'b1000110100;
    pxcRom[8683] <= 10'b1000110100;
    pxcRom[8684] <= 10'b1000110100;
    pxcRom[8685] <= 10'b1000110100;
    pxcRom[8686] <= 10'b1000110100;
    pxcRom[8687] <= 10'b1000110100;
    pxcRom[8688] <= 10'b1000110100;
    pxcRom[8689] <= 10'b1000110100;
    pxcRom[8690] <= 10'b1000000111;
    pxcRom[8691] <= 10'b1000000111;
    pxcRom[8692] <= 10'b0111101101;
    pxcRom[8693] <= 10'b0110110111;
    pxcRom[8694] <= 10'b0110000110;
    pxcRom[8695] <= 10'b0110010000;
    pxcRom[8696] <= 10'b0110001011;
    pxcRom[8697] <= 10'b0111011011;
    pxcRom[8698] <= 10'b0111101101;
    pxcRom[8699] <= 10'b1000000111;
    pxcRom[8700] <= 10'b1000000111;
    pxcRom[8701] <= 10'b1000110100;
    pxcRom[8702] <= 10'b1000110100;
    pxcRom[8703] <= 10'b1000110100;
    pxcRom[8704] <= 10'b1000110100;
    pxcRom[8705] <= 10'b1000110100;
    pxcRom[8706] <= 10'b1000110100;
    pxcRom[8707] <= 10'b1000110100;
    pxcRom[8708] <= 10'b1000110100;
    pxcRom[8709] <= 10'b1000110100;
    pxcRom[8710] <= 10'b1000000111;
    pxcRom[8711] <= 10'b1000110100;
    pxcRom[8712] <= 10'b1000110100;
    pxcRom[8713] <= 10'b1000110100;
    pxcRom[8714] <= 10'b1000110100;
    pxcRom[8715] <= 10'b1000110100;
    pxcRom[8716] <= 10'b1000110100;
    pxcRom[8717] <= 10'b0111101101;
    pxcRom[8718] <= 10'b0110110111;
    pxcRom[8719] <= 10'b0110101111;
    pxcRom[8720] <= 10'b0101100110;
    pxcRom[8721] <= 10'b0100110011;
    pxcRom[8722] <= 10'b0100011011;
    pxcRom[8723] <= 10'b0100011100;
    pxcRom[8724] <= 10'b0100100001;
    pxcRom[8725] <= 10'b0100110100;
    pxcRom[8726] <= 10'b0101000000;
    pxcRom[8727] <= 10'b0101011010;
    pxcRom[8728] <= 10'b0101111110;
    pxcRom[8729] <= 10'b0110010101;
    pxcRom[8730] <= 10'b0111000001;
    pxcRom[8731] <= 10'b0111101101;
    pxcRom[8732] <= 10'b1000110100;
    pxcRom[8733] <= 10'b1000110100;
    pxcRom[8734] <= 10'b1000110100;
    pxcRom[8735] <= 10'b1000110100;
    pxcRom[8736] <= 10'b1000110100;
    pxcRom[8737] <= 10'b1000110100;
    pxcRom[8738] <= 10'b1000000111;
    pxcRom[8739] <= 10'b1000000111;
    pxcRom[8740] <= 10'b1000000111;
    pxcRom[8741] <= 10'b0111101101;
    pxcRom[8742] <= 10'b0111011011;
    pxcRom[8743] <= 10'b0111001101;
    pxcRom[8744] <= 10'b0110011010;
    pxcRom[8745] <= 10'b0101011010;
    pxcRom[8746] <= 10'b0100010010;
    pxcRom[8747] <= 10'b0011010110;
    pxcRom[8748] <= 10'b0010011001;
    pxcRom[8749] <= 10'b0001110011;
    pxcRom[8750] <= 10'b0001011110;
    pxcRom[8751] <= 10'b0001010101;
    pxcRom[8752] <= 10'b0001010111;
    pxcRom[8753] <= 10'b0001011011;
    pxcRom[8754] <= 10'b0001100101;
    pxcRom[8755] <= 10'b0001110101;
    pxcRom[8756] <= 10'b0010001110;
    pxcRom[8757] <= 10'b0010110100;
    pxcRom[8758] <= 10'b0011101000;
    pxcRom[8759] <= 10'b0100110010;
    pxcRom[8760] <= 10'b0110000010;
    pxcRom[8761] <= 10'b1000110100;
    pxcRom[8762] <= 10'b1000110100;
    pxcRom[8763] <= 10'b1000110100;
    pxcRom[8764] <= 10'b1000110100;
    pxcRom[8765] <= 10'b1000110100;
    pxcRom[8766] <= 10'b1000000111;
    pxcRom[8767] <= 10'b0111011011;
    pxcRom[8768] <= 10'b0111011011;
    pxcRom[8769] <= 10'b0111001101;
    pxcRom[8770] <= 10'b0110100000;
    pxcRom[8771] <= 10'b0110001011;
    pxcRom[8772] <= 10'b0101110111;
    pxcRom[8773] <= 10'b0100110110;
    pxcRom[8774] <= 10'b0011110000;
    pxcRom[8775] <= 10'b0010101111;
    pxcRom[8776] <= 10'b0001111000;
    pxcRom[8777] <= 10'b0001010000;
    pxcRom[8778] <= 10'b0000111010;
    pxcRom[8779] <= 10'b0000110000;
    pxcRom[8780] <= 10'b0000101111;
    pxcRom[8781] <= 10'b0000110101;
    pxcRom[8782] <= 10'b0001000001;
    pxcRom[8783] <= 10'b0001010011;
    pxcRom[8784] <= 10'b0001101110;
    pxcRom[8785] <= 10'b0010010001;
    pxcRom[8786] <= 10'b0011001000;
    pxcRom[8787] <= 10'b0100000101;
    pxcRom[8788] <= 10'b0101011010;
    pxcRom[8789] <= 10'b1000000111;
    pxcRom[8790] <= 10'b1000000111;
    pxcRom[8791] <= 10'b1000110100;
    pxcRom[8792] <= 10'b1000110100;
    pxcRom[8793] <= 10'b1000110100;
    pxcRom[8794] <= 10'b1000110100;
    pxcRom[8795] <= 10'b0111101101;
    pxcRom[8796] <= 10'b0111011011;
    pxcRom[8797] <= 10'b0110110111;
    pxcRom[8798] <= 10'b0110100000;
    pxcRom[8799] <= 10'b0101111110;
    pxcRom[8800] <= 10'b0101010110;
    pxcRom[8801] <= 10'b0100110000;
    pxcRom[8802] <= 10'b0011101001;
    pxcRom[8803] <= 10'b0010101001;
    pxcRom[8804] <= 10'b0001110001;
    pxcRom[8805] <= 10'b0001001000;
    pxcRom[8806] <= 10'b0000110000;
    pxcRom[8807] <= 10'b0000100100;
    pxcRom[8808] <= 10'b0000100011;
    pxcRom[8809] <= 10'b0000101011;
    pxcRom[8810] <= 10'b0000111001;
    pxcRom[8811] <= 10'b0001001111;
    pxcRom[8812] <= 10'b0001101110;
    pxcRom[8813] <= 10'b0010010101;
    pxcRom[8814] <= 10'b0011001101;
    pxcRom[8815] <= 10'b0100010011;
    pxcRom[8816] <= 10'b0101011110;
    pxcRom[8817] <= 10'b1000110100;
    pxcRom[8818] <= 10'b1000110100;
    pxcRom[8819] <= 10'b1000110100;
    pxcRom[8820] <= 10'b1000110100;
    pxcRom[8821] <= 10'b1000110100;
    pxcRom[8822] <= 10'b1000000111;
    pxcRom[8823] <= 10'b0111101101;
    pxcRom[8824] <= 10'b0111001101;
    pxcRom[8825] <= 10'b0111000001;
    pxcRom[8826] <= 10'b0110101111;
    pxcRom[8827] <= 10'b0101110001;
    pxcRom[8828] <= 10'b0101010100;
    pxcRom[8829] <= 10'b0100101101;
    pxcRom[8830] <= 10'b0011110011;
    pxcRom[8831] <= 10'b0010101011;
    pxcRom[8832] <= 10'b0001101111;
    pxcRom[8833] <= 10'b0001000100;
    pxcRom[8834] <= 10'b0000101001;
    pxcRom[8835] <= 10'b0000011100;
    pxcRom[8836] <= 10'b0000011101;
    pxcRom[8837] <= 10'b0000100111;
    pxcRom[8838] <= 10'b0000111010;
    pxcRom[8839] <= 10'b0001010100;
    pxcRom[8840] <= 10'b0001111001;
    pxcRom[8841] <= 10'b0010101011;
    pxcRom[8842] <= 10'b0011100110;
    pxcRom[8843] <= 10'b0100101100;
    pxcRom[8844] <= 10'b0101110001;
    pxcRom[8845] <= 10'b1000110100;
    pxcRom[8846] <= 10'b1000000111;
    pxcRom[8847] <= 10'b1000110100;
    pxcRom[8848] <= 10'b1000110100;
    pxcRom[8849] <= 10'b1000110100;
    pxcRom[8850] <= 10'b1000110100;
    pxcRom[8851] <= 10'b1000000111;
    pxcRom[8852] <= 10'b0111011011;
    pxcRom[8853] <= 10'b0111011011;
    pxcRom[8854] <= 10'b0110000110;
    pxcRom[8855] <= 10'b0101101000;
    pxcRom[8856] <= 10'b0101010100;
    pxcRom[8857] <= 10'b0100110010;
    pxcRom[8858] <= 10'b0011111100;
    pxcRom[8859] <= 10'b0010110000;
    pxcRom[8860] <= 10'b0001101111;
    pxcRom[8861] <= 10'b0000111111;
    pxcRom[8862] <= 10'b0000100001;
    pxcRom[8863] <= 10'b0000010100;
    pxcRom[8864] <= 10'b0000010111;
    pxcRom[8865] <= 10'b0000100111;
    pxcRom[8866] <= 10'b0001000000;
    pxcRom[8867] <= 10'b0001100010;
    pxcRom[8868] <= 10'b0010010010;
    pxcRom[8869] <= 10'b0011001101;
    pxcRom[8870] <= 10'b0100001111;
    pxcRom[8871] <= 10'b0101100011;
    pxcRom[8872] <= 10'b0110100111;
    pxcRom[8873] <= 10'b1000110100;
    pxcRom[8874] <= 10'b1000110100;
    pxcRom[8875] <= 10'b1000110100;
    pxcRom[8876] <= 10'b1000110100;
    pxcRom[8877] <= 10'b1000000111;
    pxcRom[8878] <= 10'b1000110100;
    pxcRom[8879] <= 10'b1000000111;
    pxcRom[8880] <= 10'b1000000111;
    pxcRom[8881] <= 10'b0111000001;
    pxcRom[8882] <= 10'b0110000010;
    pxcRom[8883] <= 10'b0101110111;
    pxcRom[8884] <= 10'b0101011100;
    pxcRom[8885] <= 10'b0100101010;
    pxcRom[8886] <= 10'b0011111110;
    pxcRom[8887] <= 10'b0010111011;
    pxcRom[8888] <= 10'b0001110000;
    pxcRom[8889] <= 10'b0000111001;
    pxcRom[8890] <= 10'b0000011001;
    pxcRom[8891] <= 10'b0000001100;
    pxcRom[8892] <= 10'b0000010100;
    pxcRom[8893] <= 10'b0000101010;
    pxcRom[8894] <= 10'b0001001010;
    pxcRom[8895] <= 10'b0001110110;
    pxcRom[8896] <= 10'b0010110110;
    pxcRom[8897] <= 10'b0011111110;
    pxcRom[8898] <= 10'b0101001000;
    pxcRom[8899] <= 10'b0110010101;
    pxcRom[8900] <= 10'b0111000001;
    pxcRom[8901] <= 10'b1000000111;
    pxcRom[8902] <= 10'b1000000111;
    pxcRom[8903] <= 10'b1000110100;
    pxcRom[8904] <= 10'b1000110100;
    pxcRom[8905] <= 10'b1000000111;
    pxcRom[8906] <= 10'b1000110100;
    pxcRom[8907] <= 10'b1000110100;
    pxcRom[8908] <= 10'b1000000111;
    pxcRom[8909] <= 10'b0111001101;
    pxcRom[8910] <= 10'b0110100111;
    pxcRom[8911] <= 10'b0101110001;
    pxcRom[8912] <= 10'b0101011100;
    pxcRom[8913] <= 10'b0100101111;
    pxcRom[8914] <= 10'b0011111111;
    pxcRom[8915] <= 10'b0011000001;
    pxcRom[8916] <= 10'b0001101110;
    pxcRom[8917] <= 10'b0000110001;
    pxcRom[8918] <= 10'b0000001111;
    pxcRom[8919] <= 10'b0000000110;
    pxcRom[8920] <= 10'b0000010011;
    pxcRom[8921] <= 10'b0000110001;
    pxcRom[8922] <= 10'b0001011011;
    pxcRom[8923] <= 10'b0010010111;
    pxcRom[8924] <= 10'b0011101010;
    pxcRom[8925] <= 10'b0101000000;
    pxcRom[8926] <= 10'b0101110100;
    pxcRom[8927] <= 10'b0110100111;
    pxcRom[8928] <= 10'b1000110100;
    pxcRom[8929] <= 10'b0111011011;
    pxcRom[8930] <= 10'b0111101101;
    pxcRom[8931] <= 10'b1000000111;
    pxcRom[8932] <= 10'b1000110100;
    pxcRom[8933] <= 10'b1000000111;
    pxcRom[8934] <= 10'b1000000111;
    pxcRom[8935] <= 10'b1000000111;
    pxcRom[8936] <= 10'b0111001101;
    pxcRom[8937] <= 10'b0110101111;
    pxcRom[8938] <= 10'b0111000001;
    pxcRom[8939] <= 10'b0110000110;
    pxcRom[8940] <= 10'b0101101000;
    pxcRom[8941] <= 10'b0100101111;
    pxcRom[8942] <= 10'b0100000000;
    pxcRom[8943] <= 10'b0011000111;
    pxcRom[8944] <= 10'b0001101011;
    pxcRom[8945] <= 10'b0000100101;
    pxcRom[8946] <= 10'b0000000110;
    pxcRom[8947] <= 10'b0000000011;
    pxcRom[8948] <= 10'b0000010101;
    pxcRom[8949] <= 10'b0000111101;
    pxcRom[8950] <= 10'b0001111000;
    pxcRom[8951] <= 10'b0011001001;
    pxcRom[8952] <= 10'b0100101010;
    pxcRom[8953] <= 10'b0101111011;
    pxcRom[8954] <= 10'b0110010101;
    pxcRom[8955] <= 10'b0111001101;
    pxcRom[8956] <= 10'b1000000111;
    pxcRom[8957] <= 10'b0111011011;
    pxcRom[8958] <= 10'b1000000111;
    pxcRom[8959] <= 10'b1000000111;
    pxcRom[8960] <= 10'b1000110100;
    pxcRom[8961] <= 10'b1000110100;
    pxcRom[8962] <= 10'b1000110100;
    pxcRom[8963] <= 10'b1000000111;
    pxcRom[8964] <= 10'b0111001101;
    pxcRom[8965] <= 10'b0111011011;
    pxcRom[8966] <= 10'b0111000001;
    pxcRom[8967] <= 10'b0110100000;
    pxcRom[8968] <= 10'b0101010010;
    pxcRom[8969] <= 10'b0100101001;
    pxcRom[8970] <= 10'b0100000101;
    pxcRom[8971] <= 10'b0011001111;
    pxcRom[8972] <= 10'b0001100001;
    pxcRom[8973] <= 10'b0000010101;
    pxcRom[8974] <= 10'b0000000001;
    pxcRom[8975] <= 10'b0000000010;
    pxcRom[8976] <= 10'b0000011000;
    pxcRom[8977] <= 10'b0001010010;
    pxcRom[8978] <= 10'b0010100100;
    pxcRom[8979] <= 10'b0100001110;
    pxcRom[8980] <= 10'b0101110100;
    pxcRom[8981] <= 10'b0110001011;
    pxcRom[8982] <= 10'b0110110111;
    pxcRom[8983] <= 10'b0111101101;
    pxcRom[8984] <= 10'b1000110100;
    pxcRom[8985] <= 10'b1000000111;
    pxcRom[8986] <= 10'b1000110100;
    pxcRom[8987] <= 10'b1000000111;
    pxcRom[8988] <= 10'b1000110100;
    pxcRom[8989] <= 10'b1000110100;
    pxcRom[8990] <= 10'b1000110100;
    pxcRom[8991] <= 10'b0111101101;
    pxcRom[8992] <= 10'b0111011011;
    pxcRom[8993] <= 10'b0111101101;
    pxcRom[8994] <= 10'b0111001101;
    pxcRom[8995] <= 10'b0110011010;
    pxcRom[8996] <= 10'b0101011000;
    pxcRom[8997] <= 10'b0100110100;
    pxcRom[8998] <= 10'b0100010100;
    pxcRom[8999] <= 10'b0011000001;
    pxcRom[9000] <= 10'b0001001100;
    pxcRom[9001] <= 10'b0000001001;
    pxcRom[9002] <= 10'b0000000000;
    pxcRom[9003] <= 10'b0000000010;
    pxcRom[9004] <= 10'b0000100000;
    pxcRom[9005] <= 10'b0001110100;
    pxcRom[9006] <= 10'b0011100110;
    pxcRom[9007] <= 10'b0101010100;
    pxcRom[9008] <= 10'b0110010101;
    pxcRom[9009] <= 10'b0110100000;
    pxcRom[9010] <= 10'b0111001101;
    pxcRom[9011] <= 10'b1000000111;
    pxcRom[9012] <= 10'b1000110100;
    pxcRom[9013] <= 10'b1000000111;
    pxcRom[9014] <= 10'b1000110100;
    pxcRom[9015] <= 10'b1000110100;
    pxcRom[9016] <= 10'b1000110100;
    pxcRom[9017] <= 10'b1000110100;
    pxcRom[9018] <= 10'b1000110100;
    pxcRom[9019] <= 10'b0111011011;
    pxcRom[9020] <= 10'b0111011011;
    pxcRom[9021] <= 10'b0111011011;
    pxcRom[9022] <= 10'b0111001101;
    pxcRom[9023] <= 10'b0110100000;
    pxcRom[9024] <= 10'b0101011110;
    pxcRom[9025] <= 10'b0100111100;
    pxcRom[9026] <= 10'b0100001001;
    pxcRom[9027] <= 10'b0010100000;
    pxcRom[9028] <= 10'b0000110100;
    pxcRom[9029] <= 10'b0000000100;
    pxcRom[9030] <= 10'b0000000000;
    pxcRom[9031] <= 10'b0000000011;
    pxcRom[9032] <= 10'b0000110001;
    pxcRom[9033] <= 10'b0010100010;
    pxcRom[9034] <= 10'b0100100100;
    pxcRom[9035] <= 10'b0110010000;
    pxcRom[9036] <= 10'b0110100000;
    pxcRom[9037] <= 10'b0110100000;
    pxcRom[9038] <= 10'b0111000001;
    pxcRom[9039] <= 10'b1000000111;
    pxcRom[9040] <= 10'b1000000111;
    pxcRom[9041] <= 10'b1000000111;
    pxcRom[9042] <= 10'b1000110100;
    pxcRom[9043] <= 10'b1000110100;
    pxcRom[9044] <= 10'b1000110100;
    pxcRom[9045] <= 10'b1000110100;
    pxcRom[9046] <= 10'b1000000111;
    pxcRom[9047] <= 10'b0111101101;
    pxcRom[9048] <= 10'b0111011011;
    pxcRom[9049] <= 10'b1000000111;
    pxcRom[9050] <= 10'b1000000111;
    pxcRom[9051] <= 10'b0110001011;
    pxcRom[9052] <= 10'b0101101000;
    pxcRom[9053] <= 10'b0100111011;
    pxcRom[9054] <= 10'b0011011001;
    pxcRom[9055] <= 10'b0001110010;
    pxcRom[9056] <= 10'b0000100010;
    pxcRom[9057] <= 10'b0000000010;
    pxcRom[9058] <= 10'b0000000000;
    pxcRom[9059] <= 10'b0000001000;
    pxcRom[9060] <= 10'b0001001001;
    pxcRom[9061] <= 10'b0011001100;
    pxcRom[9062] <= 10'b0101010100;
    pxcRom[9063] <= 10'b0110011010;
    pxcRom[9064] <= 10'b0110110111;
    pxcRom[9065] <= 10'b0110011010;
    pxcRom[9066] <= 10'b0111000001;
    pxcRom[9067] <= 10'b1000000111;
    pxcRom[9068] <= 10'b1000000111;
    pxcRom[9069] <= 10'b1000110100;
    pxcRom[9070] <= 10'b1000110100;
    pxcRom[9071] <= 10'b1000110100;
    pxcRom[9072] <= 10'b1000110100;
    pxcRom[9073] <= 10'b1000110100;
    pxcRom[9074] <= 10'b0111101101;
    pxcRom[9075] <= 10'b1000110100;
    pxcRom[9076] <= 10'b0111101101;
    pxcRom[9077] <= 10'b0111101101;
    pxcRom[9078] <= 10'b0111000001;
    pxcRom[9079] <= 10'b0110010101;
    pxcRom[9080] <= 10'b0101011100;
    pxcRom[9081] <= 10'b0100000001;
    pxcRom[9082] <= 10'b0010011110;
    pxcRom[9083] <= 10'b0001001111;
    pxcRom[9084] <= 10'b0000011010;
    pxcRom[9085] <= 10'b0000000011;
    pxcRom[9086] <= 10'b0000000001;
    pxcRom[9087] <= 10'b0000010100;
    pxcRom[9088] <= 10'b0001011101;
    pxcRom[9089] <= 10'b0011010110;
    pxcRom[9090] <= 10'b0101010110;
    pxcRom[9091] <= 10'b0110000010;
    pxcRom[9092] <= 10'b0110010101;
    pxcRom[9093] <= 10'b0110011010;
    pxcRom[9094] <= 10'b0110101111;
    pxcRom[9095] <= 10'b0111101101;
    pxcRom[9096] <= 10'b0111011011;
    pxcRom[9097] <= 10'b1000000111;
    pxcRom[9098] <= 10'b1000000111;
    pxcRom[9099] <= 10'b1000110100;
    pxcRom[9100] <= 10'b1000110100;
    pxcRom[9101] <= 10'b1000000111;
    pxcRom[9102] <= 10'b1000000111;
    pxcRom[9103] <= 10'b1000110100;
    pxcRom[9104] <= 10'b0111101101;
    pxcRom[9105] <= 10'b0110110111;
    pxcRom[9106] <= 10'b0110100111;
    pxcRom[9107] <= 10'b0101110100;
    pxcRom[9108] <= 10'b0100010010;
    pxcRom[9109] <= 10'b0010111111;
    pxcRom[9110] <= 10'b0001110010;
    pxcRom[9111] <= 10'b0000111011;
    pxcRom[9112] <= 10'b0000010110;
    pxcRom[9113] <= 10'b0000000100;
    pxcRom[9114] <= 10'b0000000110;
    pxcRom[9115] <= 10'b0000100011;
    pxcRom[9116] <= 10'b0001101000;
    pxcRom[9117] <= 10'b0011001101;
    pxcRom[9118] <= 10'b0100101111;
    pxcRom[9119] <= 10'b0101001001;
    pxcRom[9120] <= 10'b0101110001;
    pxcRom[9121] <= 10'b0110000010;
    pxcRom[9122] <= 10'b0110000110;
    pxcRom[9123] <= 10'b0110100111;
    pxcRom[9124] <= 10'b0110101111;
    pxcRom[9125] <= 10'b0111011011;
    pxcRom[9126] <= 10'b1000000111;
    pxcRom[9127] <= 10'b1000110100;
    pxcRom[9128] <= 10'b1000110100;
    pxcRom[9129] <= 10'b1000110100;
    pxcRom[9130] <= 10'b1000110100;
    pxcRom[9131] <= 10'b1000110100;
    pxcRom[9132] <= 10'b1000110100;
    pxcRom[9133] <= 10'b0111001101;
    pxcRom[9134] <= 10'b0110000010;
    pxcRom[9135] <= 10'b0100101000;
    pxcRom[9136] <= 10'b0011011001;
    pxcRom[9137] <= 10'b0010001111;
    pxcRom[9138] <= 10'b0001011000;
    pxcRom[9139] <= 10'b0000110001;
    pxcRom[9140] <= 10'b0000010101;
    pxcRom[9141] <= 10'b0000000111;
    pxcRom[9142] <= 10'b0000001111;
    pxcRom[9143] <= 10'b0000101110;
    pxcRom[9144] <= 10'b0001101010;
    pxcRom[9145] <= 10'b0011000001;
    pxcRom[9146] <= 10'b0100001110;
    pxcRom[9147] <= 10'b0100110010;
    pxcRom[9148] <= 10'b0100111111;
    pxcRom[9149] <= 10'b0101010000;
    pxcRom[9150] <= 10'b0101110001;
    pxcRom[9151] <= 10'b0110100000;
    pxcRom[9152] <= 10'b0110101111;
    pxcRom[9153] <= 10'b0111000001;
    pxcRom[9154] <= 10'b0111101101;
    pxcRom[9155] <= 10'b0111101101;
    pxcRom[9156] <= 10'b1000110100;
    pxcRom[9157] <= 10'b1000000111;
    pxcRom[9158] <= 10'b1000000111;
    pxcRom[9159] <= 10'b0111101101;
    pxcRom[9160] <= 10'b0111101101;
    pxcRom[9161] <= 10'b0110011010;
    pxcRom[9162] <= 10'b0100110111;
    pxcRom[9163] <= 10'b0011101001;
    pxcRom[9164] <= 10'b0010100110;
    pxcRom[9165] <= 10'b0001101111;
    pxcRom[9166] <= 10'b0001000110;
    pxcRom[9167] <= 10'b0000101010;
    pxcRom[9168] <= 10'b0000010110;
    pxcRom[9169] <= 10'b0000001101;
    pxcRom[9170] <= 10'b0000011001;
    pxcRom[9171] <= 10'b0000110110;
    pxcRom[9172] <= 10'b0001100111;
    pxcRom[9173] <= 10'b0010101101;
    pxcRom[9174] <= 10'b0011110001;
    pxcRom[9175] <= 10'b0100010100;
    pxcRom[9176] <= 10'b0100110011;
    pxcRom[9177] <= 10'b0101000101;
    pxcRom[9178] <= 10'b0101101011;
    pxcRom[9179] <= 10'b0110000010;
    pxcRom[9180] <= 10'b0110100111;
    pxcRom[9181] <= 10'b0110110111;
    pxcRom[9182] <= 10'b1000000111;
    pxcRom[9183] <= 10'b0111101101;
    pxcRom[9184] <= 10'b1000110100;
    pxcRom[9185] <= 10'b1000110100;
    pxcRom[9186] <= 10'b1000110100;
    pxcRom[9187] <= 10'b0111101101;
    pxcRom[9188] <= 10'b0110110111;
    pxcRom[9189] <= 10'b0101001001;
    pxcRom[9190] <= 10'b0011110111;
    pxcRom[9191] <= 10'b0010111100;
    pxcRom[9192] <= 10'b0010000100;
    pxcRom[9193] <= 10'b0001011010;
    pxcRom[9194] <= 10'b0000111100;
    pxcRom[9195] <= 10'b0000100111;
    pxcRom[9196] <= 10'b0000011001;
    pxcRom[9197] <= 10'b0000010100;
    pxcRom[9198] <= 10'b0000100001;
    pxcRom[9199] <= 10'b0000111010;
    pxcRom[9200] <= 10'b0001100010;
    pxcRom[9201] <= 10'b0010011110;
    pxcRom[9202] <= 10'b0011011000;
    pxcRom[9203] <= 10'b0100000100;
    pxcRom[9204] <= 10'b0100100001;
    pxcRom[9205] <= 10'b0101001000;
    pxcRom[9206] <= 10'b0101101110;
    pxcRom[9207] <= 10'b0110011010;
    pxcRom[9208] <= 10'b0110100111;
    pxcRom[9209] <= 10'b0110101111;
    pxcRom[9210] <= 10'b1000000111;
    pxcRom[9211] <= 10'b1000000111;
    pxcRom[9212] <= 10'b1000110100;
    pxcRom[9213] <= 10'b1000110100;
    pxcRom[9214] <= 10'b1000000111;
    pxcRom[9215] <= 10'b0111101101;
    pxcRom[9216] <= 10'b0110000010;
    pxcRom[9217] <= 10'b0100010100;
    pxcRom[9218] <= 10'b0011010100;
    pxcRom[9219] <= 10'b0010100010;
    pxcRom[9220] <= 10'b0001110001;
    pxcRom[9221] <= 10'b0001001111;
    pxcRom[9222] <= 10'b0000110111;
    pxcRom[9223] <= 10'b0000100111;
    pxcRom[9224] <= 10'b0000011110;
    pxcRom[9225] <= 10'b0000011101;
    pxcRom[9226] <= 10'b0000100111;
    pxcRom[9227] <= 10'b0000111101;
    pxcRom[9228] <= 10'b0001011110;
    pxcRom[9229] <= 10'b0010010000;
    pxcRom[9230] <= 10'b0011001101;
    pxcRom[9231] <= 10'b0011111100;
    pxcRom[9232] <= 10'b0100100010;
    pxcRom[9233] <= 10'b0101000110;
    pxcRom[9234] <= 10'b0101111011;
    pxcRom[9235] <= 10'b0110101111;
    pxcRom[9236] <= 10'b0110110111;
    pxcRom[9237] <= 10'b0111011011;
    pxcRom[9238] <= 10'b0111101101;
    pxcRom[9239] <= 10'b1000110100;
    pxcRom[9240] <= 10'b1000110100;
    pxcRom[9241] <= 10'b1000110100;
    pxcRom[9242] <= 10'b1000000111;
    pxcRom[9243] <= 10'b0111101101;
    pxcRom[9244] <= 10'b0101101011;
    pxcRom[9245] <= 10'b0011111111;
    pxcRom[9246] <= 10'b0011000110;
    pxcRom[9247] <= 10'b0010010010;
    pxcRom[9248] <= 10'b0001100111;
    pxcRom[9249] <= 10'b0001001100;
    pxcRom[9250] <= 10'b0000110111;
    pxcRom[9251] <= 10'b0000101100;
    pxcRom[9252] <= 10'b0000100110;
    pxcRom[9253] <= 10'b0000100110;
    pxcRom[9254] <= 10'b0000101101;
    pxcRom[9255] <= 10'b0000111111;
    pxcRom[9256] <= 10'b0001011111;
    pxcRom[9257] <= 10'b0010001110;
    pxcRom[9258] <= 10'b0011001100;
    pxcRom[9259] <= 10'b0100000110;
    pxcRom[9260] <= 10'b0100111001;
    pxcRom[9261] <= 10'b0101011000;
    pxcRom[9262] <= 10'b0110101111;
    pxcRom[9263] <= 10'b0111101101;
    pxcRom[9264] <= 10'b1000000111;
    pxcRom[9265] <= 10'b0111011011;
    pxcRom[9266] <= 10'b1000000111;
    pxcRom[9267] <= 10'b1000110100;
    pxcRom[9268] <= 10'b1000110100;
    pxcRom[9269] <= 10'b1000110100;
    pxcRom[9270] <= 10'b1000110100;
    pxcRom[9271] <= 10'b1000110100;
    pxcRom[9272] <= 10'b0101100011;
    pxcRom[9273] <= 10'b0011111111;
    pxcRom[9274] <= 10'b0011001110;
    pxcRom[9275] <= 10'b0010010111;
    pxcRom[9276] <= 10'b0001101110;
    pxcRom[9277] <= 10'b0001010010;
    pxcRom[9278] <= 10'b0001000001;
    pxcRom[9279] <= 10'b0000111001;
    pxcRom[9280] <= 10'b0000110100;
    pxcRom[9281] <= 10'b0000110100;
    pxcRom[9282] <= 10'b0000111001;
    pxcRom[9283] <= 10'b0001001011;
    pxcRom[9284] <= 10'b0001101011;
    pxcRom[9285] <= 10'b0010100000;
    pxcRom[9286] <= 10'b0011100100;
    pxcRom[9287] <= 10'b0100101100;
    pxcRom[9288] <= 10'b0101100001;
    pxcRom[9289] <= 10'b0110010000;
    pxcRom[9290] <= 10'b0111001101;
    pxcRom[9291] <= 10'b1000000111;
    pxcRom[9292] <= 10'b0111011011;
    pxcRom[9293] <= 10'b1000000111;
    pxcRom[9294] <= 10'b0111011011;
    pxcRom[9295] <= 10'b1000110100;
    pxcRom[9296] <= 10'b1000110100;
    pxcRom[9297] <= 10'b1000110100;
    pxcRom[9298] <= 10'b1000110100;
    pxcRom[9299] <= 10'b1000110100;
    pxcRom[9300] <= 10'b0110100000;
    pxcRom[9301] <= 10'b0101001110;
    pxcRom[9302] <= 10'b0100010111;
    pxcRom[9303] <= 10'b0011101000;
    pxcRom[9304] <= 10'b0011000010;
    pxcRom[9305] <= 10'b0010100011;
    pxcRom[9306] <= 10'b0010010010;
    pxcRom[9307] <= 10'b0010001000;
    pxcRom[9308] <= 10'b0010000100;
    pxcRom[9309] <= 10'b0001111111;
    pxcRom[9310] <= 10'b0010000100;
    pxcRom[9311] <= 10'b0010010110;
    pxcRom[9312] <= 10'b0010111111;
    pxcRom[9313] <= 10'b0011111011;
    pxcRom[9314] <= 10'b0101001101;
    pxcRom[9315] <= 10'b0110000110;
    pxcRom[9316] <= 10'b0111011011;
    pxcRom[9317] <= 10'b0111000001;
    pxcRom[9318] <= 10'b0111101101;
    pxcRom[9319] <= 10'b0111101101;
    pxcRom[9320] <= 10'b1000110100;
    pxcRom[9321] <= 10'b1000000111;
    pxcRom[9322] <= 10'b1000110100;
    pxcRom[9323] <= 10'b1000110100;
    pxcRom[9324] <= 10'b1000110100;
    pxcRom[9325] <= 10'b1000110100;
    pxcRom[9326] <= 10'b1000110100;
    pxcRom[9327] <= 10'b1000110100;
    pxcRom[9328] <= 10'b1000110100;
    pxcRom[9329] <= 10'b1000000111;
    pxcRom[9330] <= 10'b1000000111;
    pxcRom[9331] <= 10'b0110110111;
    pxcRom[9332] <= 10'b0110100000;
    pxcRom[9333] <= 10'b0110001011;
    pxcRom[9334] <= 10'b0110000110;
    pxcRom[9335] <= 10'b0101101110;
    pxcRom[9336] <= 10'b0101010110;
    pxcRom[9337] <= 10'b0101001000;
    pxcRom[9338] <= 10'b0101001001;
    pxcRom[9339] <= 10'b0101111011;
    pxcRom[9340] <= 10'b0110100000;
    pxcRom[9341] <= 10'b0111101101;
    pxcRom[9342] <= 10'b1000110100;
    pxcRom[9343] <= 10'b1000110100;
    pxcRom[9344] <= 10'b1000110100;
    pxcRom[9345] <= 10'b1000110100;
    pxcRom[9346] <= 10'b1000110100;
    pxcRom[9347] <= 10'b1000110100;
    pxcRom[9348] <= 10'b1000110100;
    pxcRom[9349] <= 10'b1000110100;
    pxcRom[9350] <= 10'b1000110100;
    pxcRom[9351] <= 10'b1000110100;
    pxcRom[9352] <= 10'b1000110100;
    pxcRom[9353] <= 10'b1000110100;
    pxcRom[9354] <= 10'b1000110100;
    pxcRom[9355] <= 10'b1000110100;
    pxcRom[9356] <= 10'b1000110100;
    pxcRom[9357] <= 10'b1000110100;
    pxcRom[9358] <= 10'b1000110100;
    pxcRom[9359] <= 10'b1000110100;
    pxcRom[9360] <= 10'b1000110100;
    pxcRom[9361] <= 10'b1000110100;
    pxcRom[9362] <= 10'b1000000111;
    pxcRom[9363] <= 10'b1000000111;
    pxcRom[9364] <= 10'b1000110100;
    pxcRom[9365] <= 10'b1000110100;
    pxcRom[9366] <= 10'b1000000111;
    pxcRom[9367] <= 10'b1000000111;
    pxcRom[9368] <= 10'b1000000111;
    pxcRom[9369] <= 10'b1000110100;
    pxcRom[9370] <= 10'b1000110100;
    pxcRom[9371] <= 10'b1000110100;
    pxcRom[9372] <= 10'b1000110100;
    pxcRom[9373] <= 10'b1000110100;
    pxcRom[9374] <= 10'b1000110100;
    pxcRom[9375] <= 10'b1000110100;
    pxcRom[9376] <= 10'b1000110100;
    pxcRom[9377] <= 10'b1000110100;
    pxcRom[9378] <= 10'b1000110100;
    pxcRom[9379] <= 10'b1000110100;
    pxcRom[9380] <= 10'b1000110100;
    pxcRom[9381] <= 10'b1000110100;
    pxcRom[9382] <= 10'b1000110100;
    pxcRom[9383] <= 10'b1000110100;
    pxcRom[9384] <= 10'b1000110100;
    pxcRom[9385] <= 10'b1000110100;
    pxcRom[9386] <= 10'b1000110100;
    pxcRom[9387] <= 10'b1000110100;
    pxcRom[9388] <= 10'b1000110100;
    pxcRom[9389] <= 10'b1000110100;
    pxcRom[9390] <= 10'b1000110100;
    pxcRom[9391] <= 10'b1000110100;
    pxcRom[9392] <= 10'b1000110100;
    pxcRom[9393] <= 10'b1000110100;
    pxcRom[9394] <= 10'b1000110100;
    pxcRom[9395] <= 10'b1000110100;
    pxcRom[9396] <= 10'b1000110100;
    pxcRom[9397] <= 10'b1000110100;
    pxcRom[9398] <= 10'b1000110100;
    pxcRom[9399] <= 10'b1000110100;
    pxcRom[9400] <= 10'b1000110100;
    pxcRom[9401] <= 10'b1000110100;
    pxcRom[9402] <= 10'b1000110100;
    pxcRom[9403] <= 10'b1000110100;
    pxcRom[9404] <= 10'b1000110100;
    pxcRom[9405] <= 10'b1000110100;
    pxcRom[9406] <= 10'b1000110100;
    pxcRom[9407] <= 10'b1000110100;
    pxcRom[9408] <= 10'b1000101100;
    pxcRom[9409] <= 10'b1000101100;
    pxcRom[9410] <= 10'b1000101100;
    pxcRom[9411] <= 10'b1000101100;
    pxcRom[9412] <= 10'b1000101100;
    pxcRom[9413] <= 10'b1000101100;
    pxcRom[9414] <= 10'b1000101100;
    pxcRom[9415] <= 10'b1000101100;
    pxcRom[9416] <= 10'b1000101100;
    pxcRom[9417] <= 10'b1000101100;
    pxcRom[9418] <= 10'b1000101100;
    pxcRom[9419] <= 10'b1000101100;
    pxcRom[9420] <= 10'b1000101100;
    pxcRom[9421] <= 10'b0111111111;
    pxcRom[9422] <= 10'b0111111111;
    pxcRom[9423] <= 10'b1000101100;
    pxcRom[9424] <= 10'b1000101100;
    pxcRom[9425] <= 10'b1000101100;
    pxcRom[9426] <= 10'b1000101100;
    pxcRom[9427] <= 10'b1000101100;
    pxcRom[9428] <= 10'b1000101100;
    pxcRom[9429] <= 10'b1000101100;
    pxcRom[9430] <= 10'b1000101100;
    pxcRom[9431] <= 10'b1000101100;
    pxcRom[9432] <= 10'b1000101100;
    pxcRom[9433] <= 10'b1000101100;
    pxcRom[9434] <= 10'b1000101100;
    pxcRom[9435] <= 10'b1000101100;
    pxcRom[9436] <= 10'b1000101100;
    pxcRom[9437] <= 10'b1000101100;
    pxcRom[9438] <= 10'b1000101100;
    pxcRom[9439] <= 10'b1000101100;
    pxcRom[9440] <= 10'b1000101100;
    pxcRom[9441] <= 10'b1000101100;
    pxcRom[9442] <= 10'b1000101100;
    pxcRom[9443] <= 10'b1000101100;
    pxcRom[9444] <= 10'b0111100110;
    pxcRom[9445] <= 10'b0111010011;
    pxcRom[9446] <= 10'b0110111001;
    pxcRom[9447] <= 10'b0111000101;
    pxcRom[9448] <= 10'b0111010011;
    pxcRom[9449] <= 10'b0110111001;
    pxcRom[9450] <= 10'b0110101111;
    pxcRom[9451] <= 10'b0110011000;
    pxcRom[9452] <= 10'b0110001101;
    pxcRom[9453] <= 10'b0110101111;
    pxcRom[9454] <= 10'b0111111111;
    pxcRom[9455] <= 10'b1000101100;
    pxcRom[9456] <= 10'b1000101100;
    pxcRom[9457] <= 10'b1000101100;
    pxcRom[9458] <= 10'b1000101100;
    pxcRom[9459] <= 10'b1000101100;
    pxcRom[9460] <= 10'b1000101100;
    pxcRom[9461] <= 10'b1000101100;
    pxcRom[9462] <= 10'b1000101100;
    pxcRom[9463] <= 10'b1000101100;
    pxcRom[9464] <= 10'b1000101100;
    pxcRom[9465] <= 10'b1000101100;
    pxcRom[9466] <= 10'b1000101100;
    pxcRom[9467] <= 10'b1000101100;
    pxcRom[9468] <= 10'b1000101100;
    pxcRom[9469] <= 10'b0111111111;
    pxcRom[9470] <= 10'b0111000101;
    pxcRom[9471] <= 10'b0110010010;
    pxcRom[9472] <= 10'b0101100110;
    pxcRom[9473] <= 10'b0100111000;
    pxcRom[9474] <= 10'b0100100010;
    pxcRom[9475] <= 10'b0100001010;
    pxcRom[9476] <= 10'b0011111000;
    pxcRom[9477] <= 10'b0011110100;
    pxcRom[9478] <= 10'b0011101101;
    pxcRom[9479] <= 10'b0011110000;
    pxcRom[9480] <= 10'b0011111101;
    pxcRom[9481] <= 10'b0100011000;
    pxcRom[9482] <= 10'b0100111000;
    pxcRom[9483] <= 10'b0101101111;
    pxcRom[9484] <= 10'b0110100111;
    pxcRom[9485] <= 10'b0111100110;
    pxcRom[9486] <= 10'b1000101100;
    pxcRom[9487] <= 10'b0111111111;
    pxcRom[9488] <= 10'b0111100110;
    pxcRom[9489] <= 10'b0111111111;
    pxcRom[9490] <= 10'b1000101100;
    pxcRom[9491] <= 10'b1000101100;
    pxcRom[9492] <= 10'b1000101100;
    pxcRom[9493] <= 10'b1000101100;
    pxcRom[9494] <= 10'b1000101100;
    pxcRom[9495] <= 10'b1000101100;
    pxcRom[9496] <= 10'b0111111111;
    pxcRom[9497] <= 10'b0101111010;
    pxcRom[9498] <= 10'b0100110011;
    pxcRom[9499] <= 10'b0011111100;
    pxcRom[9500] <= 10'b0011001110;
    pxcRom[9501] <= 10'b0010101000;
    pxcRom[9502] <= 10'b0010010000;
    pxcRom[9503] <= 10'b0001111010;
    pxcRom[9504] <= 10'b0001101011;
    pxcRom[9505] <= 10'b0001100001;
    pxcRom[9506] <= 10'b0001011100;
    pxcRom[9507] <= 10'b0001011110;
    pxcRom[9508] <= 10'b0001100101;
    pxcRom[9509] <= 10'b0001110101;
    pxcRom[9510] <= 10'b0010001101;
    pxcRom[9511] <= 10'b0010101101;
    pxcRom[9512] <= 10'b0011010000;
    pxcRom[9513] <= 10'b0100000011;
    pxcRom[9514] <= 10'b0101001100;
    pxcRom[9515] <= 10'b0110111001;
    pxcRom[9516] <= 10'b0111100110;
    pxcRom[9517] <= 10'b0111111111;
    pxcRom[9518] <= 10'b1000101100;
    pxcRom[9519] <= 10'b1000101100;
    pxcRom[9520] <= 10'b1000101100;
    pxcRom[9521] <= 10'b1000101100;
    pxcRom[9522] <= 10'b0111111111;
    pxcRom[9523] <= 10'b0111100110;
    pxcRom[9524] <= 10'b0110010010;
    pxcRom[9525] <= 10'b0100011101;
    pxcRom[9526] <= 10'b0011011100;
    pxcRom[9527] <= 10'b0010101010;
    pxcRom[9528] <= 10'b0010000011;
    pxcRom[9529] <= 10'b0001100011;
    pxcRom[9530] <= 10'b0001001101;
    pxcRom[9531] <= 10'b0000111010;
    pxcRom[9532] <= 10'b0000101101;
    pxcRom[9533] <= 10'b0000100100;
    pxcRom[9534] <= 10'b0000100001;
    pxcRom[9535] <= 10'b0000100010;
    pxcRom[9536] <= 10'b0000100111;
    pxcRom[9537] <= 10'b0000110010;
    pxcRom[9538] <= 10'b0001000101;
    pxcRom[9539] <= 10'b0001011111;
    pxcRom[9540] <= 10'b0010000001;
    pxcRom[9541] <= 10'b0010101110;
    pxcRom[9542] <= 10'b0011101100;
    pxcRom[9543] <= 10'b0101011110;
    pxcRom[9544] <= 10'b0111100110;
    pxcRom[9545] <= 10'b0111100110;
    pxcRom[9546] <= 10'b1000101100;
    pxcRom[9547] <= 10'b1000101100;
    pxcRom[9548] <= 10'b1000101100;
    pxcRom[9549] <= 10'b1000101100;
    pxcRom[9550] <= 10'b0111100110;
    pxcRom[9551] <= 10'b0111010011;
    pxcRom[9552] <= 10'b0101000110;
    pxcRom[9553] <= 10'b0011100110;
    pxcRom[9554] <= 10'b0010100111;
    pxcRom[9555] <= 10'b0001111011;
    pxcRom[9556] <= 10'b0001011010;
    pxcRom[9557] <= 10'b0001000010;
    pxcRom[9558] <= 10'b0000101111;
    pxcRom[9559] <= 10'b0000100010;
    pxcRom[9560] <= 10'b0000011001;
    pxcRom[9561] <= 10'b0000010011;
    pxcRom[9562] <= 10'b0000010001;
    pxcRom[9563] <= 10'b0000010000;
    pxcRom[9564] <= 10'b0000010100;
    pxcRom[9565] <= 10'b0000011011;
    pxcRom[9566] <= 10'b0000101010;
    pxcRom[9567] <= 10'b0000111111;
    pxcRom[9568] <= 10'b0001011100;
    pxcRom[9569] <= 10'b0010000001;
    pxcRom[9570] <= 10'b0010110111;
    pxcRom[9571] <= 10'b0100011000;
    pxcRom[9572] <= 10'b0110101111;
    pxcRom[9573] <= 10'b0111100110;
    pxcRom[9574] <= 10'b1000101100;
    pxcRom[9575] <= 10'b1000101100;
    pxcRom[9576] <= 10'b1000101100;
    pxcRom[9577] <= 10'b1000101100;
    pxcRom[9578] <= 10'b0111111111;
    pxcRom[9579] <= 10'b0110011111;
    pxcRom[9580] <= 10'b0100100000;
    pxcRom[9581] <= 10'b0011000101;
    pxcRom[9582] <= 10'b0010001000;
    pxcRom[9583] <= 10'b0001100011;
    pxcRom[9584] <= 10'b0001000111;
    pxcRom[9585] <= 10'b0000110100;
    pxcRom[9586] <= 10'b0000100101;
    pxcRom[9587] <= 10'b0000011100;
    pxcRom[9588] <= 10'b0000010110;
    pxcRom[9589] <= 10'b0000010011;
    pxcRom[9590] <= 10'b0000010001;
    pxcRom[9591] <= 10'b0000010000;
    pxcRom[9592] <= 10'b0000010001;
    pxcRom[9593] <= 10'b0000010101;
    pxcRom[9594] <= 10'b0000011110;
    pxcRom[9595] <= 10'b0000101111;
    pxcRom[9596] <= 10'b0001001000;
    pxcRom[9597] <= 10'b0001101001;
    pxcRom[9598] <= 10'b0010011101;
    pxcRom[9599] <= 10'b0011110100;
    pxcRom[9600] <= 10'b0110101111;
    pxcRom[9601] <= 10'b0111111111;
    pxcRom[9602] <= 10'b0111111111;
    pxcRom[9603] <= 10'b1000101100;
    pxcRom[9604] <= 10'b1000101100;
    pxcRom[9605] <= 10'b1000101100;
    pxcRom[9606] <= 10'b0111100110;
    pxcRom[9607] <= 10'b0110001000;
    pxcRom[9608] <= 10'b0100000110;
    pxcRom[9609] <= 10'b0010110010;
    pxcRom[9610] <= 10'b0001111011;
    pxcRom[9611] <= 10'b0001011010;
    pxcRom[9612] <= 10'b0001000011;
    pxcRom[9613] <= 10'b0000110011;
    pxcRom[9614] <= 10'b0000101000;
    pxcRom[9615] <= 10'b0000100010;
    pxcRom[9616] <= 10'b0000100000;
    pxcRom[9617] <= 10'b0000100000;
    pxcRom[9618] <= 10'b0000011111;
    pxcRom[9619] <= 10'b0000011101;
    pxcRom[9620] <= 10'b0000011001;
    pxcRom[9621] <= 10'b0000011000;
    pxcRom[9622] <= 10'b0000011100;
    pxcRom[9623] <= 10'b0000101000;
    pxcRom[9624] <= 10'b0000111110;
    pxcRom[9625] <= 10'b0001011100;
    pxcRom[9626] <= 10'b0010001001;
    pxcRom[9627] <= 10'b0011011110;
    pxcRom[9628] <= 10'b0110011000;
    pxcRom[9629] <= 10'b0111100110;
    pxcRom[9630] <= 10'b0111111111;
    pxcRom[9631] <= 10'b1000101100;
    pxcRom[9632] <= 10'b1000101100;
    pxcRom[9633] <= 10'b0111111111;
    pxcRom[9634] <= 10'b0111010011;
    pxcRom[9635] <= 10'b0110001101;
    pxcRom[9636] <= 10'b0100000011;
    pxcRom[9637] <= 10'b0010101100;
    pxcRom[9638] <= 10'b0001111011;
    pxcRom[9639] <= 10'b0001011110;
    pxcRom[9640] <= 10'b0001001100;
    pxcRom[9641] <= 10'b0000111110;
    pxcRom[9642] <= 10'b0000110110;
    pxcRom[9643] <= 10'b0000110101;
    pxcRom[9644] <= 10'b0000110101;
    pxcRom[9645] <= 10'b0000110110;
    pxcRom[9646] <= 10'b0000110100;
    pxcRom[9647] <= 10'b0000101111;
    pxcRom[9648] <= 10'b0000100101;
    pxcRom[9649] <= 10'b0000011101;
    pxcRom[9650] <= 10'b0000011100;
    pxcRom[9651] <= 10'b0000100100;
    pxcRom[9652] <= 10'b0000111000;
    pxcRom[9653] <= 10'b0001010110;
    pxcRom[9654] <= 10'b0010000011;
    pxcRom[9655] <= 10'b0011011001;
    pxcRom[9656] <= 10'b0110011111;
    pxcRom[9657] <= 10'b0111010011;
    pxcRom[9658] <= 10'b1000101100;
    pxcRom[9659] <= 10'b1000101100;
    pxcRom[9660] <= 10'b1000101100;
    pxcRom[9661] <= 10'b1000101100;
    pxcRom[9662] <= 10'b0111010011;
    pxcRom[9663] <= 10'b0101111111;
    pxcRom[9664] <= 10'b0100000000;
    pxcRom[9665] <= 10'b0010110011;
    pxcRom[9666] <= 10'b0010000100;
    pxcRom[9667] <= 10'b0001101110;
    pxcRom[9668] <= 10'b0001011110;
    pxcRom[9669] <= 10'b0001010100;
    pxcRom[9670] <= 10'b0001001110;
    pxcRom[9671] <= 10'b0001010000;
    pxcRom[9672] <= 10'b0001010011;
    pxcRom[9673] <= 10'b0001010101;
    pxcRom[9674] <= 10'b0001001111;
    pxcRom[9675] <= 10'b0001000000;
    pxcRom[9676] <= 10'b0000101101;
    pxcRom[9677] <= 10'b0000100000;
    pxcRom[9678] <= 10'b0000011011;
    pxcRom[9679] <= 10'b0000100011;
    pxcRom[9680] <= 10'b0000110110;
    pxcRom[9681] <= 10'b0001010111;
    pxcRom[9682] <= 10'b0010000010;
    pxcRom[9683] <= 10'b0011010101;
    pxcRom[9684] <= 10'b0110101111;
    pxcRom[9685] <= 10'b0111111111;
    pxcRom[9686] <= 10'b0111111111;
    pxcRom[9687] <= 10'b1000101100;
    pxcRom[9688] <= 10'b1000101100;
    pxcRom[9689] <= 10'b1000101100;
    pxcRom[9690] <= 10'b0111100110;
    pxcRom[9691] <= 10'b0110001101;
    pxcRom[9692] <= 10'b0100011011;
    pxcRom[9693] <= 10'b0011000100;
    pxcRom[9694] <= 10'b0010011100;
    pxcRom[9695] <= 10'b0010000111;
    pxcRom[9696] <= 10'b0001111000;
    pxcRom[9697] <= 10'b0001110001;
    pxcRom[9698] <= 10'b0001110000;
    pxcRom[9699] <= 10'b0001110011;
    pxcRom[9700] <= 10'b0001110111;
    pxcRom[9701] <= 10'b0001110111;
    pxcRom[9702] <= 10'b0001100011;
    pxcRom[9703] <= 10'b0001001000;
    pxcRom[9704] <= 10'b0000101111;
    pxcRom[9705] <= 10'b0000011111;
    pxcRom[9706] <= 10'b0000011011;
    pxcRom[9707] <= 10'b0000100011;
    pxcRom[9708] <= 10'b0000111000;
    pxcRom[9709] <= 10'b0001011010;
    pxcRom[9710] <= 10'b0010001010;
    pxcRom[9711] <= 10'b0011011101;
    pxcRom[9712] <= 10'b0101111010;
    pxcRom[9713] <= 10'b0110111001;
    pxcRom[9714] <= 10'b0111010011;
    pxcRom[9715] <= 10'b1000101100;
    pxcRom[9716] <= 10'b1000101100;
    pxcRom[9717] <= 10'b1000101100;
    pxcRom[9718] <= 10'b1000101100;
    pxcRom[9719] <= 10'b0110100111;
    pxcRom[9720] <= 10'b0100110000;
    pxcRom[9721] <= 10'b0011100001;
    pxcRom[9722] <= 10'b0010111100;
    pxcRom[9723] <= 10'b0010101100;
    pxcRom[9724] <= 10'b0010011110;
    pxcRom[9725] <= 10'b0010010110;
    pxcRom[9726] <= 10'b0010010011;
    pxcRom[9727] <= 10'b0010010111;
    pxcRom[9728] <= 10'b0010010100;
    pxcRom[9729] <= 10'b0010000101;
    pxcRom[9730] <= 10'b0001100100;
    pxcRom[9731] <= 10'b0001000011;
    pxcRom[9732] <= 10'b0000101010;
    pxcRom[9733] <= 10'b0000011101;
    pxcRom[9734] <= 10'b0000011011;
    pxcRom[9735] <= 10'b0000100101;
    pxcRom[9736] <= 10'b0000111101;
    pxcRom[9737] <= 10'b0001100010;
    pxcRom[9738] <= 10'b0010011000;
    pxcRom[9739] <= 10'b0011101001;
    pxcRom[9740] <= 10'b0101001100;
    pxcRom[9741] <= 10'b0101111010;
    pxcRom[9742] <= 10'b0111010011;
    pxcRom[9743] <= 10'b1000101100;
    pxcRom[9744] <= 10'b1000101100;
    pxcRom[9745] <= 10'b1000101100;
    pxcRom[9746] <= 10'b1000101100;
    pxcRom[9747] <= 10'b0111000101;
    pxcRom[9748] <= 10'b0101010100;
    pxcRom[9749] <= 10'b0100000111;
    pxcRom[9750] <= 10'b0011101001;
    pxcRom[9751] <= 10'b0011001110;
    pxcRom[9752] <= 10'b0010111011;
    pxcRom[9753] <= 10'b0010101111;
    pxcRom[9754] <= 10'b0010100100;
    pxcRom[9755] <= 10'b0010011001;
    pxcRom[9756] <= 10'b0010001011;
    pxcRom[9757] <= 10'b0001101110;
    pxcRom[9758] <= 10'b0001001111;
    pxcRom[9759] <= 10'b0000110110;
    pxcRom[9760] <= 10'b0000100100;
    pxcRom[9761] <= 10'b0000011011;
    pxcRom[9762] <= 10'b0000011100;
    pxcRom[9763] <= 10'b0000101010;
    pxcRom[9764] <= 10'b0001000101;
    pxcRom[9765] <= 10'b0001101111;
    pxcRom[9766] <= 10'b0010100111;
    pxcRom[9767] <= 10'b0011110111;
    pxcRom[9768] <= 10'b0100101010;
    pxcRom[9769] <= 10'b0101010010;
    pxcRom[9770] <= 10'b0110101111;
    pxcRom[9771] <= 10'b0111111111;
    pxcRom[9772] <= 10'b1000101100;
    pxcRom[9773] <= 10'b1000101100;
    pxcRom[9774] <= 10'b0111111111;
    pxcRom[9775] <= 10'b0111010011;
    pxcRom[9776] <= 10'b0101100011;
    pxcRom[9777] <= 10'b0100011000;
    pxcRom[9778] <= 10'b0011100101;
    pxcRom[9779] <= 10'b0011000001;
    pxcRom[9780] <= 10'b0010100111;
    pxcRom[9781] <= 10'b0010010010;
    pxcRom[9782] <= 10'b0001111111;
    pxcRom[9783] <= 10'b0001101101;
    pxcRom[9784] <= 10'b0001011100;
    pxcRom[9785] <= 10'b0001001001;
    pxcRom[9786] <= 10'b0000110111;
    pxcRom[9787] <= 10'b0000101000;
    pxcRom[9788] <= 10'b0000011101;
    pxcRom[9789] <= 10'b0000011001;
    pxcRom[9790] <= 10'b0000100001;
    pxcRom[9791] <= 10'b0000110011;
    pxcRom[9792] <= 10'b0001010000;
    pxcRom[9793] <= 10'b0001111110;
    pxcRom[9794] <= 10'b0010110100;
    pxcRom[9795] <= 10'b0011101001;
    pxcRom[9796] <= 10'b0100000101;
    pxcRom[9797] <= 10'b0100100110;
    pxcRom[9798] <= 10'b0101100110;
    pxcRom[9799] <= 10'b0111010011;
    pxcRom[9800] <= 10'b1000101100;
    pxcRom[9801] <= 10'b1000101100;
    pxcRom[9802] <= 10'b1000101100;
    pxcRom[9803] <= 10'b0110100111;
    pxcRom[9804] <= 10'b0100111101;
    pxcRom[9805] <= 10'b0011101010;
    pxcRom[9806] <= 10'b0010110100;
    pxcRom[9807] <= 10'b0010001111;
    pxcRom[9808] <= 10'b0001110100;
    pxcRom[9809] <= 10'b0001100000;
    pxcRom[9810] <= 10'b0001001111;
    pxcRom[9811] <= 10'b0001000000;
    pxcRom[9812] <= 10'b0000110100;
    pxcRom[9813] <= 10'b0000101001;
    pxcRom[9814] <= 10'b0000100000;
    pxcRom[9815] <= 10'b0000011001;
    pxcRom[9816] <= 10'b0000010111;
    pxcRom[9817] <= 10'b0000011010;
    pxcRom[9818] <= 10'b0000100101;
    pxcRom[9819] <= 10'b0000111010;
    pxcRom[9820] <= 10'b0001011100;
    pxcRom[9821] <= 10'b0010000110;
    pxcRom[9822] <= 10'b0010110001;
    pxcRom[9823] <= 10'b0011010000;
    pxcRom[9824] <= 10'b0011100101;
    pxcRom[9825] <= 10'b0100000110;
    pxcRom[9826] <= 10'b0101000110;
    pxcRom[9827] <= 10'b0111100110;
    pxcRom[9828] <= 10'b1000101100;
    pxcRom[9829] <= 10'b1000101100;
    pxcRom[9830] <= 10'b0111111111;
    pxcRom[9831] <= 10'b0101100000;
    pxcRom[9832] <= 10'b0011110111;
    pxcRom[9833] <= 10'b0010101111;
    pxcRom[9834] <= 10'b0001111111;
    pxcRom[9835] <= 10'b0001100000;
    pxcRom[9836] <= 10'b0001001010;
    pxcRom[9837] <= 10'b0000111011;
    pxcRom[9838] <= 10'b0000101110;
    pxcRom[9839] <= 10'b0000100100;
    pxcRom[9840] <= 10'b0000011011;
    pxcRom[9841] <= 10'b0000010100;
    pxcRom[9842] <= 10'b0000010001;
    pxcRom[9843] <= 10'b0000010000;
    pxcRom[9844] <= 10'b0000010100;
    pxcRom[9845] <= 10'b0000011100;
    pxcRom[9846] <= 10'b0000101011;
    pxcRom[9847] <= 10'b0001000000;
    pxcRom[9848] <= 10'b0001011101;
    pxcRom[9849] <= 10'b0001111011;
    pxcRom[9850] <= 10'b0010010111;
    pxcRom[9851] <= 10'b0010101010;
    pxcRom[9852] <= 10'b0011000001;
    pxcRom[9853] <= 10'b0011101011;
    pxcRom[9854] <= 10'b0100110001;
    pxcRom[9855] <= 10'b0110101111;
    pxcRom[9856] <= 10'b1000101100;
    pxcRom[9857] <= 10'b1000101100;
    pxcRom[9858] <= 10'b0111000101;
    pxcRom[9859] <= 10'b0100100010;
    pxcRom[9860] <= 10'b0010111111;
    pxcRom[9861] <= 10'b0010000000;
    pxcRom[9862] <= 10'b0001011010;
    pxcRom[9863] <= 10'b0001000001;
    pxcRom[9864] <= 10'b0000110000;
    pxcRom[9865] <= 10'b0000100100;
    pxcRom[9866] <= 10'b0000011100;
    pxcRom[9867] <= 10'b0000010110;
    pxcRom[9868] <= 10'b0000010000;
    pxcRom[9869] <= 10'b0000001101;
    pxcRom[9870] <= 10'b0000001100;
    pxcRom[9871] <= 10'b0000001111;
    pxcRom[9872] <= 10'b0000010101;
    pxcRom[9873] <= 10'b0000011111;
    pxcRom[9874] <= 10'b0000101100;
    pxcRom[9875] <= 10'b0000111111;
    pxcRom[9876] <= 10'b0001010011;
    pxcRom[9877] <= 10'b0001100111;
    pxcRom[9878] <= 10'b0001110111;
    pxcRom[9879] <= 10'b0010000111;
    pxcRom[9880] <= 10'b0010011111;
    pxcRom[9881] <= 10'b0011000111;
    pxcRom[9882] <= 10'b0100011010;
    pxcRom[9883] <= 10'b0110111001;
    pxcRom[9884] <= 10'b1000101100;
    pxcRom[9885] <= 10'b1000101100;
    pxcRom[9886] <= 10'b0110111001;
    pxcRom[9887] <= 10'b0011101110;
    pxcRom[9888] <= 10'b0010011000;
    pxcRom[9889] <= 10'b0001100010;
    pxcRom[9890] <= 10'b0001000010;
    pxcRom[9891] <= 10'b0000101110;
    pxcRom[9892] <= 10'b0000100100;
    pxcRom[9893] <= 10'b0000011100;
    pxcRom[9894] <= 10'b0000010111;
    pxcRom[9895] <= 10'b0000010010;
    pxcRom[9896] <= 10'b0000001111;
    pxcRom[9897] <= 10'b0000001101;
    pxcRom[9898] <= 10'b0000001110;
    pxcRom[9899] <= 10'b0000010001;
    pxcRom[9900] <= 10'b0000010111;
    pxcRom[9901] <= 10'b0000011111;
    pxcRom[9902] <= 10'b0000101000;
    pxcRom[9903] <= 10'b0000110101;
    pxcRom[9904] <= 10'b0001000001;
    pxcRom[9905] <= 10'b0001001110;
    pxcRom[9906] <= 10'b0001011011;
    pxcRom[9907] <= 10'b0001101101;
    pxcRom[9908] <= 10'b0010000100;
    pxcRom[9909] <= 10'b0010101111;
    pxcRom[9910] <= 10'b0100010100;
    pxcRom[9911] <= 10'b0110111001;
    pxcRom[9912] <= 10'b1000101100;
    pxcRom[9913] <= 10'b1000101100;
    pxcRom[9914] <= 10'b0110011111;
    pxcRom[9915] <= 10'b0011001111;
    pxcRom[9916] <= 10'b0010000000;
    pxcRom[9917] <= 10'b0001010010;
    pxcRom[9918] <= 10'b0000110101;
    pxcRom[9919] <= 10'b0000100101;
    pxcRom[9920] <= 10'b0000011101;
    pxcRom[9921] <= 10'b0000011000;
    pxcRom[9922] <= 10'b0000010100;
    pxcRom[9923] <= 10'b0000010010;
    pxcRom[9924] <= 10'b0000001111;
    pxcRom[9925] <= 10'b0000001111;
    pxcRom[9926] <= 10'b0000010000;
    pxcRom[9927] <= 10'b0000010011;
    pxcRom[9928] <= 10'b0000010111;
    pxcRom[9929] <= 10'b0000011011;
    pxcRom[9930] <= 10'b0000100001;
    pxcRom[9931] <= 10'b0000101001;
    pxcRom[9932] <= 10'b0000110001;
    pxcRom[9933] <= 10'b0000111011;
    pxcRom[9934] <= 10'b0001000111;
    pxcRom[9935] <= 10'b0001011000;
    pxcRom[9936] <= 10'b0001110011;
    pxcRom[9937] <= 10'b0010101000;
    pxcRom[9938] <= 10'b0100100010;
    pxcRom[9939] <= 10'b0111000101;
    pxcRom[9940] <= 10'b1000101100;
    pxcRom[9941] <= 10'b1000101100;
    pxcRom[9942] <= 10'b0110010010;
    pxcRom[9943] <= 10'b0011000000;
    pxcRom[9944] <= 10'b0001110100;
    pxcRom[9945] <= 10'b0001001011;
    pxcRom[9946] <= 10'b0000101111;
    pxcRom[9947] <= 10'b0000011111;
    pxcRom[9948] <= 10'b0000010110;
    pxcRom[9949] <= 10'b0000010010;
    pxcRom[9950] <= 10'b0000001111;
    pxcRom[9951] <= 10'b0000001110;
    pxcRom[9952] <= 10'b0000001110;
    pxcRom[9953] <= 10'b0000010000;
    pxcRom[9954] <= 10'b0000010010;
    pxcRom[9955] <= 10'b0000010110;
    pxcRom[9956] <= 10'b0000011001;
    pxcRom[9957] <= 10'b0000011100;
    pxcRom[9958] <= 10'b0000011110;
    pxcRom[9959] <= 10'b0000100010;
    pxcRom[9960] <= 10'b0000101001;
    pxcRom[9961] <= 10'b0000110001;
    pxcRom[9962] <= 10'b0000111111;
    pxcRom[9963] <= 10'b0001010011;
    pxcRom[9964] <= 10'b0001110010;
    pxcRom[9965] <= 10'b0010101111;
    pxcRom[9966] <= 10'b0100101010;
    pxcRom[9967] <= 10'b0111100110;
    pxcRom[9968] <= 10'b1000101100;
    pxcRom[9969] <= 10'b1000101100;
    pxcRom[9970] <= 10'b0101101111;
    pxcRom[9971] <= 10'b0010111100;
    pxcRom[9972] <= 10'b0001110101;
    pxcRom[9973] <= 10'b0001001100;
    pxcRom[9974] <= 10'b0000101111;
    pxcRom[9975] <= 10'b0000011110;
    pxcRom[9976] <= 10'b0000010011;
    pxcRom[9977] <= 10'b0000001110;
    pxcRom[9978] <= 10'b0000001101;
    pxcRom[9979] <= 10'b0000001101;
    pxcRom[9980] <= 10'b0000010000;
    pxcRom[9981] <= 10'b0000010101;
    pxcRom[9982] <= 10'b0000011011;
    pxcRom[9983] <= 10'b0000011111;
    pxcRom[9984] <= 10'b0000100001;
    pxcRom[9985] <= 10'b0000100010;
    pxcRom[9986] <= 10'b0000100011;
    pxcRom[9987] <= 10'b0000100101;
    pxcRom[9988] <= 10'b0000101010;
    pxcRom[9989] <= 10'b0000110100;
    pxcRom[9990] <= 10'b0001000011;
    pxcRom[9991] <= 10'b0001011011;
    pxcRom[9992] <= 10'b0001111111;
    pxcRom[9993] <= 10'b0011000011;
    pxcRom[9994] <= 10'b0100111011;
    pxcRom[9995] <= 10'b1000101100;
    pxcRom[9996] <= 10'b1000101100;
    pxcRom[9997] <= 10'b0111111111;
    pxcRom[9998] <= 10'b0101101111;
    pxcRom[9999] <= 10'b0011001011;
    pxcRom[10000] <= 10'b0010000001;
    pxcRom[10001] <= 10'b0001010111;
    pxcRom[10002] <= 10'b0000111001;
    pxcRom[10003] <= 10'b0000100101;
    pxcRom[10004] <= 10'b0000011001;
    pxcRom[10005] <= 10'b0000010011;
    pxcRom[10006] <= 10'b0000010010;
    pxcRom[10007] <= 10'b0000010101;
    pxcRom[10008] <= 10'b0000011011;
    pxcRom[10009] <= 10'b0000100010;
    pxcRom[10010] <= 10'b0000101011;
    pxcRom[10011] <= 10'b0000110001;
    pxcRom[10012] <= 10'b0000110100;
    pxcRom[10013] <= 10'b0000110011;
    pxcRom[10014] <= 10'b0000110010;
    pxcRom[10015] <= 10'b0000110010;
    pxcRom[10016] <= 10'b0000111000;
    pxcRom[10017] <= 10'b0001000100;
    pxcRom[10018] <= 10'b0001010111;
    pxcRom[10019] <= 10'b0001110000;
    pxcRom[10020] <= 10'b0010011001;
    pxcRom[10021] <= 10'b0011100111;
    pxcRom[10022] <= 10'b0101101100;
    pxcRom[10023] <= 10'b1000101100;
    pxcRom[10024] <= 10'b1000101100;
    pxcRom[10025] <= 10'b1000101100;
    pxcRom[10026] <= 10'b0110001101;
    pxcRom[10027] <= 10'b0011110000;
    pxcRom[10028] <= 10'b0010100010;
    pxcRom[10029] <= 10'b0001110101;
    pxcRom[10030] <= 10'b0001010001;
    pxcRom[10031] <= 10'b0000111011;
    pxcRom[10032] <= 10'b0000101101;
    pxcRom[10033] <= 10'b0000100111;
    pxcRom[10034] <= 10'b0000100110;
    pxcRom[10035] <= 10'b0000101011;
    pxcRom[10036] <= 10'b0000110011;
    pxcRom[10037] <= 10'b0000111110;
    pxcRom[10038] <= 10'b0001001000;
    pxcRom[10039] <= 10'b0001001111;
    pxcRom[10040] <= 10'b0001010001;
    pxcRom[10041] <= 10'b0001001111;
    pxcRom[10042] <= 10'b0001001110;
    pxcRom[10043] <= 10'b0001010000;
    pxcRom[10044] <= 10'b0001010110;
    pxcRom[10045] <= 10'b0001100100;
    pxcRom[10046] <= 10'b0001111000;
    pxcRom[10047] <= 10'b0010010110;
    pxcRom[10048] <= 10'b0011000100;
    pxcRom[10049] <= 10'b0100010101;
    pxcRom[10050] <= 10'b0111010011;
    pxcRom[10051] <= 10'b1000101100;
    pxcRom[10052] <= 10'b1000101100;
    pxcRom[10053] <= 10'b1000101100;
    pxcRom[10054] <= 10'b0111111111;
    pxcRom[10055] <= 10'b0101001010;
    pxcRom[10056] <= 10'b0011110000;
    pxcRom[10057] <= 10'b0010111000;
    pxcRom[10058] <= 10'b0010010010;
    pxcRom[10059] <= 10'b0001110111;
    pxcRom[10060] <= 10'b0001100111;
    pxcRom[10061] <= 10'b0001011110;
    pxcRom[10062] <= 10'b0001011101;
    pxcRom[10063] <= 10'b0001100010;
    pxcRom[10064] <= 10'b0001101010;
    pxcRom[10065] <= 10'b0001110110;
    pxcRom[10066] <= 10'b0001111111;
    pxcRom[10067] <= 10'b0010000111;
    pxcRom[10068] <= 10'b0010001000;
    pxcRom[10069] <= 10'b0010001000;
    pxcRom[10070] <= 10'b0010001000;
    pxcRom[10071] <= 10'b0010001100;
    pxcRom[10072] <= 10'b0010010010;
    pxcRom[10073] <= 10'b0010100000;
    pxcRom[10074] <= 10'b0010110111;
    pxcRom[10075] <= 10'b0011011000;
    pxcRom[10076] <= 10'b0100011110;
    pxcRom[10077] <= 10'b0110001000;
    pxcRom[10078] <= 10'b0111111111;
    pxcRom[10079] <= 10'b1000101100;
    pxcRom[10080] <= 10'b1000101100;
    pxcRom[10081] <= 10'b1000101100;
    pxcRom[10082] <= 10'b1000101100;
    pxcRom[10083] <= 10'b0111111111;
    pxcRom[10084] <= 10'b0110010010;
    pxcRom[10085] <= 10'b0101011011;
    pxcRom[10086] <= 10'b0100101110;
    pxcRom[10087] <= 10'b0100010000;
    pxcRom[10088] <= 10'b0011111110;
    pxcRom[10089] <= 10'b0011110101;
    pxcRom[10090] <= 10'b0011101011;
    pxcRom[10091] <= 10'b0011101010;
    pxcRom[10092] <= 10'b0011100101;
    pxcRom[10093] <= 10'b0011101011;
    pxcRom[10094] <= 10'b0011101011;
    pxcRom[10095] <= 10'b0011101110;
    pxcRom[10096] <= 10'b0011110000;
    pxcRom[10097] <= 10'b0011110001;
    pxcRom[10098] <= 10'b0011111001;
    pxcRom[10099] <= 10'b0100000100;
    pxcRom[10100] <= 10'b0100010001;
    pxcRom[10101] <= 10'b0100011101;
    pxcRom[10102] <= 10'b0100101111;
    pxcRom[10103] <= 10'b0101000011;
    pxcRom[10104] <= 10'b0101111010;
    pxcRom[10105] <= 10'b0110111001;
    pxcRom[10106] <= 10'b0111111111;
    pxcRom[10107] <= 10'b1000101100;
    pxcRom[10108] <= 10'b1000101100;
    pxcRom[10109] <= 10'b1000101100;
    pxcRom[10110] <= 10'b1000101100;
    pxcRom[10111] <= 10'b1000101100;
    pxcRom[10112] <= 10'b1000101100;
    pxcRom[10113] <= 10'b1000101100;
    pxcRom[10114] <= 10'b0111111111;
    pxcRom[10115] <= 10'b0111100110;
    pxcRom[10116] <= 10'b0111100110;
    pxcRom[10117] <= 10'b0111100110;
    pxcRom[10118] <= 10'b0111000101;
    pxcRom[10119] <= 10'b0110101111;
    pxcRom[10120] <= 10'b0110011111;
    pxcRom[10121] <= 10'b0110001000;
    pxcRom[10122] <= 10'b0101111010;
    pxcRom[10123] <= 10'b0101110111;
    pxcRom[10124] <= 10'b0101111111;
    pxcRom[10125] <= 10'b0101111010;
    pxcRom[10126] <= 10'b0110001000;
    pxcRom[10127] <= 10'b0110011000;
    pxcRom[10128] <= 10'b0110100111;
    pxcRom[10129] <= 10'b0110111001;
    pxcRom[10130] <= 10'b0111010011;
    pxcRom[10131] <= 10'b0111111111;
    pxcRom[10132] <= 10'b1000101100;
    pxcRom[10133] <= 10'b0111111111;
    pxcRom[10134] <= 10'b0111111111;
    pxcRom[10135] <= 10'b1000101100;
    pxcRom[10136] <= 10'b1000101100;
    pxcRom[10137] <= 10'b1000101100;
    pxcRom[10138] <= 10'b1000101100;
    pxcRom[10139] <= 10'b1000101100;
    pxcRom[10140] <= 10'b1000101100;
    pxcRom[10141] <= 10'b1000101100;
    pxcRom[10142] <= 10'b1000101100;
    pxcRom[10143] <= 10'b1000101100;
    pxcRom[10144] <= 10'b1000101100;
    pxcRom[10145] <= 10'b1000101100;
    pxcRom[10146] <= 10'b1000101100;
    pxcRom[10147] <= 10'b1000101100;
    pxcRom[10148] <= 10'b1000101100;
    pxcRom[10149] <= 10'b1000101100;
    pxcRom[10150] <= 10'b1000101100;
    pxcRom[10151] <= 10'b1000101100;
    pxcRom[10152] <= 10'b1000101100;
    pxcRom[10153] <= 10'b1000101100;
    pxcRom[10154] <= 10'b1000101100;
    pxcRom[10155] <= 10'b1000101100;
    pxcRom[10156] <= 10'b1000101100;
    pxcRom[10157] <= 10'b1000101100;
    pxcRom[10158] <= 10'b1000101100;
    pxcRom[10159] <= 10'b1000101100;
    pxcRom[10160] <= 10'b1000101100;
    pxcRom[10161] <= 10'b1000101100;
    pxcRom[10162] <= 10'b1000101100;
    pxcRom[10163] <= 10'b1000101100;
    pxcRom[10164] <= 10'b1000101100;
    pxcRom[10165] <= 10'b1000101100;
    pxcRom[10166] <= 10'b1000101100;
    pxcRom[10167] <= 10'b1000101100;
    pxcRom[10168] <= 10'b1000101100;
    pxcRom[10169] <= 10'b1000101100;
    pxcRom[10170] <= 10'b1000101100;
    pxcRom[10171] <= 10'b1000101100;
    pxcRom[10172] <= 10'b1000101100;
    pxcRom[10173] <= 10'b1000101100;
    pxcRom[10174] <= 10'b1000101100;
    pxcRom[10175] <= 10'b1000101100;
    pxcRom[10176] <= 10'b1000101100;
    pxcRom[10177] <= 10'b1000101100;
    pxcRom[10178] <= 10'b1000101100;
    pxcRom[10179] <= 10'b1000101100;
    pxcRom[10180] <= 10'b1000101100;
    pxcRom[10181] <= 10'b1000101100;
    pxcRom[10182] <= 10'b1000101100;
    pxcRom[10183] <= 10'b1000101100;
    pxcRom[10184] <= 10'b1000101100;
    pxcRom[10185] <= 10'b1000101100;
    pxcRom[10186] <= 10'b1000101100;
    pxcRom[10187] <= 10'b1000101100;
    pxcRom[10188] <= 10'b1000101100;
    pxcRom[10189] <= 10'b1000101100;
    pxcRom[10190] <= 10'b1000101100;
    pxcRom[10191] <= 10'b1000101100;
    pxcRom[10192] <= 10'b1000101110;
    pxcRom[10193] <= 10'b1000101110;
    pxcRom[10194] <= 10'b1000101110;
    pxcRom[10195] <= 10'b1000101110;
    pxcRom[10196] <= 10'b1000101110;
    pxcRom[10197] <= 10'b1000101110;
    pxcRom[10198] <= 10'b1000101110;
    pxcRom[10199] <= 10'b1000101110;
    pxcRom[10200] <= 10'b1000101110;
    pxcRom[10201] <= 10'b1000101110;
    pxcRom[10202] <= 10'b1000101110;
    pxcRom[10203] <= 10'b1000101110;
    pxcRom[10204] <= 10'b1000101110;
    pxcRom[10205] <= 10'b1000101110;
    pxcRom[10206] <= 10'b1000101110;
    pxcRom[10207] <= 10'b1000101110;
    pxcRom[10208] <= 10'b1000101110;
    pxcRom[10209] <= 10'b1000101110;
    pxcRom[10210] <= 10'b1000101110;
    pxcRom[10211] <= 10'b1000101110;
    pxcRom[10212] <= 10'b1000101110;
    pxcRom[10213] <= 10'b1000101110;
    pxcRom[10214] <= 10'b1000101110;
    pxcRom[10215] <= 10'b1000101110;
    pxcRom[10216] <= 10'b1000101110;
    pxcRom[10217] <= 10'b1000101110;
    pxcRom[10218] <= 10'b1000101110;
    pxcRom[10219] <= 10'b1000101110;
    pxcRom[10220] <= 10'b1000101110;
    pxcRom[10221] <= 10'b1000101110;
    pxcRom[10222] <= 10'b1000101110;
    pxcRom[10223] <= 10'b1000101110;
    pxcRom[10224] <= 10'b1000101110;
    pxcRom[10225] <= 10'b1000101110;
    pxcRom[10226] <= 10'b1000101110;
    pxcRom[10227] <= 10'b1000101110;
    pxcRom[10228] <= 10'b1000101110;
    pxcRom[10229] <= 10'b1000101110;
    pxcRom[10230] <= 10'b1000101110;
    pxcRom[10231] <= 10'b1000101110;
    pxcRom[10232] <= 10'b1000101110;
    pxcRom[10233] <= 10'b1000101110;
    pxcRom[10234] <= 10'b1000101110;
    pxcRom[10235] <= 10'b1000101110;
    pxcRom[10236] <= 10'b1000101110;
    pxcRom[10237] <= 10'b1000101110;
    pxcRom[10238] <= 10'b1000101110;
    pxcRom[10239] <= 10'b1000101110;
    pxcRom[10240] <= 10'b1000101110;
    pxcRom[10241] <= 10'b1000101110;
    pxcRom[10242] <= 10'b1000101110;
    pxcRom[10243] <= 10'b1000101110;
    pxcRom[10244] <= 10'b1000101110;
    pxcRom[10245] <= 10'b1000101110;
    pxcRom[10246] <= 10'b1000101110;
    pxcRom[10247] <= 10'b1000101110;
    pxcRom[10248] <= 10'b1000101110;
    pxcRom[10249] <= 10'b1000101110;
    pxcRom[10250] <= 10'b1000101110;
    pxcRom[10251] <= 10'b1000101110;
    pxcRom[10252] <= 10'b1000101110;
    pxcRom[10253] <= 10'b1000101110;
    pxcRom[10254] <= 10'b1000101110;
    pxcRom[10255] <= 10'b1000101110;
    pxcRom[10256] <= 10'b1000101110;
    pxcRom[10257] <= 10'b1000101110;
    pxcRom[10258] <= 10'b1000000001;
    pxcRom[10259] <= 10'b0111100111;
    pxcRom[10260] <= 10'b0111100111;
    pxcRom[10261] <= 10'b0111100111;
    pxcRom[10262] <= 10'b0111100111;
    pxcRom[10263] <= 10'b0111010101;
    pxcRom[10264] <= 10'b0111100111;
    pxcRom[10265] <= 10'b0111100111;
    pxcRom[10266] <= 10'b0111100111;
    pxcRom[10267] <= 10'b1000000001;
    pxcRom[10268] <= 10'b1000101110;
    pxcRom[10269] <= 10'b1000101110;
    pxcRom[10270] <= 10'b1000101110;
    pxcRom[10271] <= 10'b1000101110;
    pxcRom[10272] <= 10'b1000101110;
    pxcRom[10273] <= 10'b1000101110;
    pxcRom[10274] <= 10'b1000101110;
    pxcRom[10275] <= 10'b1000101110;
    pxcRom[10276] <= 10'b1000101110;
    pxcRom[10277] <= 10'b1000101110;
    pxcRom[10278] <= 10'b1000101110;
    pxcRom[10279] <= 10'b1000101110;
    pxcRom[10280] <= 10'b1000101110;
    pxcRom[10281] <= 10'b0110111011;
    pxcRom[10282] <= 10'b0110101001;
    pxcRom[10283] <= 10'b0110000000;
    pxcRom[10284] <= 10'b0101001010;
    pxcRom[10285] <= 10'b0100101001;
    pxcRom[10286] <= 10'b0100001100;
    pxcRom[10287] <= 10'b0011101110;
    pxcRom[10288] <= 10'b0011011110;
    pxcRom[10289] <= 10'b0011010110;
    pxcRom[10290] <= 10'b0011010010;
    pxcRom[10291] <= 10'b0011010100;
    pxcRom[10292] <= 10'b0011011110;
    pxcRom[10293] <= 10'b0011101001;
    pxcRom[10294] <= 10'b0011111101;
    pxcRom[10295] <= 10'b0100100101;
    pxcRom[10296] <= 10'b0101000000;
    pxcRom[10297] <= 10'b0101110001;
    pxcRom[10298] <= 10'b0111000111;
    pxcRom[10299] <= 10'b1000101110;
    pxcRom[10300] <= 10'b1000101110;
    pxcRom[10301] <= 10'b1000101110;
    pxcRom[10302] <= 10'b1000101110;
    pxcRom[10303] <= 10'b1000101110;
    pxcRom[10304] <= 10'b1000101110;
    pxcRom[10305] <= 10'b1000000001;
    pxcRom[10306] <= 10'b1000000001;
    pxcRom[10307] <= 10'b0111000111;
    pxcRom[10308] <= 10'b0101111100;
    pxcRom[10309] <= 10'b0100011110;
    pxcRom[10310] <= 10'b0011101011;
    pxcRom[10311] <= 10'b0010111111;
    pxcRom[10312] <= 10'b0010011010;
    pxcRom[10313] <= 10'b0001111100;
    pxcRom[10314] <= 10'b0001100110;
    pxcRom[10315] <= 10'b0001010110;
    pxcRom[10316] <= 10'b0001001100;
    pxcRom[10317] <= 10'b0001000101;
    pxcRom[10318] <= 10'b0001000100;
    pxcRom[10319] <= 10'b0001000111;
    pxcRom[10320] <= 10'b0001010001;
    pxcRom[10321] <= 10'b0001100001;
    pxcRom[10322] <= 10'b0001110111;
    pxcRom[10323] <= 10'b0010010010;
    pxcRom[10324] <= 10'b0010111001;
    pxcRom[10325] <= 10'b0011101101;
    pxcRom[10326] <= 10'b0100101011;
    pxcRom[10327] <= 10'b0110101001;
    pxcRom[10328] <= 10'b1000101110;
    pxcRom[10329] <= 10'b1000101110;
    pxcRom[10330] <= 10'b1000101110;
    pxcRom[10331] <= 10'b1000101110;
    pxcRom[10332] <= 10'b1000101110;
    pxcRom[10333] <= 10'b1000101110;
    pxcRom[10334] <= 10'b1000000001;
    pxcRom[10335] <= 10'b0101110101;
    pxcRom[10336] <= 10'b0100000001;
    pxcRom[10337] <= 10'b0011000011;
    pxcRom[10338] <= 10'b0010010101;
    pxcRom[10339] <= 10'b0001110000;
    pxcRom[10340] <= 10'b0001010011;
    pxcRom[10341] <= 10'b0000111011;
    pxcRom[10342] <= 10'b0000101010;
    pxcRom[10343] <= 10'b0000011110;
    pxcRom[10344] <= 10'b0000010110;
    pxcRom[10345] <= 10'b0000010001;
    pxcRom[10346] <= 10'b0000010001;
    pxcRom[10347] <= 10'b0000010011;
    pxcRom[10348] <= 10'b0000011001;
    pxcRom[10349] <= 10'b0000100101;
    pxcRom[10350] <= 10'b0000111000;
    pxcRom[10351] <= 10'b0001010000;
    pxcRom[10352] <= 10'b0001101111;
    pxcRom[10353] <= 10'b0010011010;
    pxcRom[10354] <= 10'b0011011111;
    pxcRom[10355] <= 10'b0101000010;
    pxcRom[10356] <= 10'b0110111011;
    pxcRom[10357] <= 10'b1000101110;
    pxcRom[10358] <= 10'b1000101110;
    pxcRom[10359] <= 10'b1000101110;
    pxcRom[10360] <= 10'b1000101110;
    pxcRom[10361] <= 10'b1000101110;
    pxcRom[10362] <= 10'b0110110001;
    pxcRom[10363] <= 10'b0100100010;
    pxcRom[10364] <= 10'b0011001100;
    pxcRom[10365] <= 10'b0010010110;
    pxcRom[10366] <= 10'b0001101111;
    pxcRom[10367] <= 10'b0001001111;
    pxcRom[10368] <= 10'b0000110110;
    pxcRom[10369] <= 10'b0000100100;
    pxcRom[10370] <= 10'b0000011000;
    pxcRom[10371] <= 10'b0000010001;
    pxcRom[10372] <= 10'b0000001100;
    pxcRom[10373] <= 10'b0000001001;
    pxcRom[10374] <= 10'b0000001000;
    pxcRom[10375] <= 10'b0000001000;
    pxcRom[10376] <= 10'b0000001011;
    pxcRom[10377] <= 10'b0000010011;
    pxcRom[10378] <= 10'b0000100001;
    pxcRom[10379] <= 10'b0000110101;
    pxcRom[10380] <= 10'b0001010000;
    pxcRom[10381] <= 10'b0001110110;
    pxcRom[10382] <= 10'b0010110010;
    pxcRom[10383] <= 10'b0100010001;
    pxcRom[10384] <= 10'b0110011010;
    pxcRom[10385] <= 10'b1000101110;
    pxcRom[10386] <= 10'b1000101110;
    pxcRom[10387] <= 10'b1000101110;
    pxcRom[10388] <= 10'b1000101110;
    pxcRom[10389] <= 10'b0111000111;
    pxcRom[10390] <= 10'b0110110001;
    pxcRom[10391] <= 10'b0100000001;
    pxcRom[10392] <= 10'b0010110100;
    pxcRom[10393] <= 10'b0010000110;
    pxcRom[10394] <= 10'b0001100010;
    pxcRom[10395] <= 10'b0001001000;
    pxcRom[10396] <= 10'b0000110100;
    pxcRom[10397] <= 10'b0000100110;
    pxcRom[10398] <= 10'b0000011110;
    pxcRom[10399] <= 10'b0000011001;
    pxcRom[10400] <= 10'b0000010111;
    pxcRom[10401] <= 10'b0000010110;
    pxcRom[10402] <= 10'b0000010011;
    pxcRom[10403] <= 10'b0000001111;
    pxcRom[10404] <= 10'b0000001110;
    pxcRom[10405] <= 10'b0000010001;
    pxcRom[10406] <= 10'b0000011011;
    pxcRom[10407] <= 10'b0000101011;
    pxcRom[10408] <= 10'b0001000100;
    pxcRom[10409] <= 10'b0001100110;
    pxcRom[10410] <= 10'b0010011111;
    pxcRom[10411] <= 10'b0011111101;
    pxcRom[10412] <= 10'b0110010100;
    pxcRom[10413] <= 10'b1000101110;
    pxcRom[10414] <= 10'b1000101110;
    pxcRom[10415] <= 10'b1000101110;
    pxcRom[10416] <= 10'b1000101110;
    pxcRom[10417] <= 10'b1000000001;
    pxcRom[10418] <= 10'b0110110001;
    pxcRom[10419] <= 10'b0011110111;
    pxcRom[10420] <= 10'b0010110100;
    pxcRom[10421] <= 10'b0010001011;
    pxcRom[10422] <= 10'b0001101010;
    pxcRom[10423] <= 10'b0001010100;
    pxcRom[10424] <= 10'b0001000100;
    pxcRom[10425] <= 10'b0000111001;
    pxcRom[10426] <= 10'b0000110110;
    pxcRom[10427] <= 10'b0000110101;
    pxcRom[10428] <= 10'b0000110110;
    pxcRom[10429] <= 10'b0000110100;
    pxcRom[10430] <= 10'b0000101011;
    pxcRom[10431] <= 10'b0000011111;
    pxcRom[10432] <= 10'b0000011000;
    pxcRom[10433] <= 10'b0000010101;
    pxcRom[10434] <= 10'b0000011010;
    pxcRom[10435] <= 10'b0000101001;
    pxcRom[10436] <= 10'b0001000010;
    pxcRom[10437] <= 10'b0001100101;
    pxcRom[10438] <= 10'b0010011101;
    pxcRom[10439] <= 10'b0011111011;
    pxcRom[10440] <= 10'b0110101001;
    pxcRom[10441] <= 10'b1000101110;
    pxcRom[10442] <= 10'b1000101110;
    pxcRom[10443] <= 10'b1000101110;
    pxcRom[10444] <= 10'b1000101110;
    pxcRom[10445] <= 10'b1000000001;
    pxcRom[10446] <= 10'b0110101001;
    pxcRom[10447] <= 10'b0100001010;
    pxcRom[10448] <= 10'b0011000011;
    pxcRom[10449] <= 10'b0010100000;
    pxcRom[10450] <= 10'b0010000000;
    pxcRom[10451] <= 10'b0001101111;
    pxcRom[10452] <= 10'b0001100100;
    pxcRom[10453] <= 10'b0001011101;
    pxcRom[10454] <= 10'b0001011100;
    pxcRom[10455] <= 10'b0001011011;
    pxcRom[10456] <= 10'b0001010111;
    pxcRom[10457] <= 10'b0001001011;
    pxcRom[10458] <= 10'b0000111000;
    pxcRom[10459] <= 10'b0000100101;
    pxcRom[10460] <= 10'b0000011000;
    pxcRom[10461] <= 10'b0000010101;
    pxcRom[10462] <= 10'b0000011100;
    pxcRom[10463] <= 10'b0000101101;
    pxcRom[10464] <= 10'b0001001000;
    pxcRom[10465] <= 10'b0001110010;
    pxcRom[10466] <= 10'b0010101011;
    pxcRom[10467] <= 10'b0100001011;
    pxcRom[10468] <= 10'b0111010101;
    pxcRom[10469] <= 10'b1000000001;
    pxcRom[10470] <= 10'b1000101110;
    pxcRom[10471] <= 10'b1000101110;
    pxcRom[10472] <= 10'b1000101110;
    pxcRom[10473] <= 10'b1000000001;
    pxcRom[10474] <= 10'b0110111011;
    pxcRom[10475] <= 10'b0100100001;
    pxcRom[10476] <= 10'b0011100111;
    pxcRom[10477] <= 10'b0011000110;
    pxcRom[10478] <= 10'b0010101010;
    pxcRom[10479] <= 10'b0010011011;
    pxcRom[10480] <= 10'b0010001101;
    pxcRom[10481] <= 10'b0010000101;
    pxcRom[10482] <= 10'b0001111000;
    pxcRom[10483] <= 10'b0001100111;
    pxcRom[10484] <= 10'b0001010010;
    pxcRom[10485] <= 10'b0000111100;
    pxcRom[10486] <= 10'b0000100110;
    pxcRom[10487] <= 10'b0000011000;
    pxcRom[10488] <= 10'b0000010001;
    pxcRom[10489] <= 10'b0000010100;
    pxcRom[10490] <= 10'b0000100000;
    pxcRom[10491] <= 10'b0000110111;
    pxcRom[10492] <= 10'b0001011001;
    pxcRom[10493] <= 10'b0010001010;
    pxcRom[10494] <= 10'b0011000110;
    pxcRom[10495] <= 10'b0100110011;
    pxcRom[10496] <= 10'b1000000001;
    pxcRom[10497] <= 10'b0111100111;
    pxcRom[10498] <= 10'b1000101110;
    pxcRom[10499] <= 10'b1000101110;
    pxcRom[10500] <= 10'b1000101110;
    pxcRom[10501] <= 10'b1000000001;
    pxcRom[10502] <= 10'b0111000111;
    pxcRom[10503] <= 10'b0101000111;
    pxcRom[10504] <= 10'b0100001110;
    pxcRom[10505] <= 10'b0011110011;
    pxcRom[10506] <= 10'b0011011000;
    pxcRom[10507] <= 10'b0010111111;
    pxcRom[10508] <= 10'b0010100100;
    pxcRom[10509] <= 10'b0010000011;
    pxcRom[10510] <= 10'b0001100010;
    pxcRom[10511] <= 10'b0001000010;
    pxcRom[10512] <= 10'b0000101101;
    pxcRom[10513] <= 10'b0000011100;
    pxcRom[10514] <= 10'b0000010010;
    pxcRom[10515] <= 10'b0000001100;
    pxcRom[10516] <= 10'b0000001101;
    pxcRom[10517] <= 10'b0000010101;
    pxcRom[10518] <= 10'b0000100111;
    pxcRom[10519] <= 10'b0001000110;
    pxcRom[10520] <= 10'b0001101110;
    pxcRom[10521] <= 10'b0010101001;
    pxcRom[10522] <= 10'b0011111111;
    pxcRom[10523] <= 10'b0101100010;
    pxcRom[10524] <= 10'b1000101110;
    pxcRom[10525] <= 10'b1000000001;
    pxcRom[10526] <= 10'b1000101110;
    pxcRom[10527] <= 10'b1000101110;
    pxcRom[10528] <= 10'b1000101110;
    pxcRom[10529] <= 10'b1000101110;
    pxcRom[10530] <= 10'b1000101110;
    pxcRom[10531] <= 10'b0101111100;
    pxcRom[10532] <= 10'b0100110111;
    pxcRom[10533] <= 10'b0100010000;
    pxcRom[10534] <= 10'b0011110110;
    pxcRom[10535] <= 10'b0011000011;
    pxcRom[10536] <= 10'b0010001101;
    pxcRom[10537] <= 10'b0001011110;
    pxcRom[10538] <= 10'b0000111011;
    pxcRom[10539] <= 10'b0000100011;
    pxcRom[10540] <= 10'b0000010100;
    pxcRom[10541] <= 10'b0000001011;
    pxcRom[10542] <= 10'b0000000111;
    pxcRom[10543] <= 10'b0000000111;
    pxcRom[10544] <= 10'b0000001011;
    pxcRom[10545] <= 10'b0000010101;
    pxcRom[10546] <= 10'b0000101011;
    pxcRom[10547] <= 10'b0001001010;
    pxcRom[10548] <= 10'b0001111001;
    pxcRom[10549] <= 10'b0010111001;
    pxcRom[10550] <= 10'b0100001000;
    pxcRom[10551] <= 10'b0110000000;
    pxcRom[10552] <= 10'b1000000001;
    pxcRom[10553] <= 10'b0111100111;
    pxcRom[10554] <= 10'b1000101110;
    pxcRom[10555] <= 10'b1000101110;
    pxcRom[10556] <= 10'b1000101110;
    pxcRom[10557] <= 10'b1000101110;
    pxcRom[10558] <= 10'b1000101110;
    pxcRom[10559] <= 10'b0110110001;
    pxcRom[10560] <= 10'b0101011011;
    pxcRom[10561] <= 10'b0100110000;
    pxcRom[10562] <= 10'b0011110000;
    pxcRom[10563] <= 10'b0010101100;
    pxcRom[10564] <= 10'b0001110110;
    pxcRom[10565] <= 10'b0001001000;
    pxcRom[10566] <= 10'b0000101001;
    pxcRom[10567] <= 10'b0000010110;
    pxcRom[10568] <= 10'b0000001100;
    pxcRom[10569] <= 10'b0000001000;
    pxcRom[10570] <= 10'b0000000111;
    pxcRom[10571] <= 10'b0000001000;
    pxcRom[10572] <= 10'b0000001100;
    pxcRom[10573] <= 10'b0000010100;
    pxcRom[10574] <= 10'b0000100100;
    pxcRom[10575] <= 10'b0000111110;
    pxcRom[10576] <= 10'b0001100111;
    pxcRom[10577] <= 10'b0010011110;
    pxcRom[10578] <= 10'b0011101100;
    pxcRom[10579] <= 10'b0101001110;
    pxcRom[10580] <= 10'b0111010101;
    pxcRom[10581] <= 10'b1000000001;
    pxcRom[10582] <= 10'b1000101110;
    pxcRom[10583] <= 10'b1000101110;
    pxcRom[10584] <= 10'b1000101110;
    pxcRom[10585] <= 10'b0111100111;
    pxcRom[10586] <= 10'b1000000001;
    pxcRom[10587] <= 10'b0110100001;
    pxcRom[10588] <= 10'b0101001110;
    pxcRom[10589] <= 10'b0100011100;
    pxcRom[10590] <= 10'b0011100011;
    pxcRom[10591] <= 10'b0010100100;
    pxcRom[10592] <= 10'b0001101110;
    pxcRom[10593] <= 10'b0001000110;
    pxcRom[10594] <= 10'b0000101011;
    pxcRom[10595] <= 10'b0000011011;
    pxcRom[10596] <= 10'b0000010011;
    pxcRom[10597] <= 10'b0000010001;
    pxcRom[10598] <= 10'b0000010001;
    pxcRom[10599] <= 10'b0000010010;
    pxcRom[10600] <= 10'b0000010001;
    pxcRom[10601] <= 10'b0000010011;
    pxcRom[10602] <= 10'b0000011010;
    pxcRom[10603] <= 10'b0000101101;
    pxcRom[10604] <= 10'b0001001101;
    pxcRom[10605] <= 10'b0001111101;
    pxcRom[10606] <= 10'b0010111010;
    pxcRom[10607] <= 10'b0100010110;
    pxcRom[10608] <= 10'b0110011010;
    pxcRom[10609] <= 10'b1000000001;
    pxcRom[10610] <= 10'b1000101110;
    pxcRom[10611] <= 10'b1000101110;
    pxcRom[10612] <= 10'b1000101110;
    pxcRom[10613] <= 10'b1000000001;
    pxcRom[10614] <= 10'b0110011010;
    pxcRom[10615] <= 10'b0101010010;
    pxcRom[10616] <= 10'b0100100110;
    pxcRom[10617] <= 10'b0011111011;
    pxcRom[10618] <= 10'b0011010110;
    pxcRom[10619] <= 10'b0010101100;
    pxcRom[10620] <= 10'b0001111100;
    pxcRom[10621] <= 10'b0001010110;
    pxcRom[10622] <= 10'b0000111110;
    pxcRom[10623] <= 10'b0000110001;
    pxcRom[10624] <= 10'b0000101100;
    pxcRom[10625] <= 10'b0000101011;
    pxcRom[10626] <= 10'b0000101010;
    pxcRom[10627] <= 10'b0000100110;
    pxcRom[10628] <= 10'b0000011111;
    pxcRom[10629] <= 10'b0000010111;
    pxcRom[10630] <= 10'b0000010111;
    pxcRom[10631] <= 10'b0000100001;
    pxcRom[10632] <= 10'b0000111001;
    pxcRom[10633] <= 10'b0001100011;
    pxcRom[10634] <= 10'b0010010111;
    pxcRom[10635] <= 10'b0011100101;
    pxcRom[10636] <= 10'b0101101011;
    pxcRom[10637] <= 10'b1000101110;
    pxcRom[10638] <= 10'b0111100111;
    pxcRom[10639] <= 10'b1000101110;
    pxcRom[10640] <= 10'b1000101110;
    pxcRom[10641] <= 10'b0111100111;
    pxcRom[10642] <= 10'b0101100000;
    pxcRom[10643] <= 10'b0100010111;
    pxcRom[10644] <= 10'b0011101110;
    pxcRom[10645] <= 10'b0011010101;
    pxcRom[10646] <= 10'b0011000100;
    pxcRom[10647] <= 10'b0010110000;
    pxcRom[10648] <= 10'b0010010010;
    pxcRom[10649] <= 10'b0001110111;
    pxcRom[10650] <= 10'b0001100101;
    pxcRom[10651] <= 10'b0001011010;
    pxcRom[10652] <= 10'b0001011000;
    pxcRom[10653] <= 10'b0001011000;
    pxcRom[10654] <= 10'b0001010010;
    pxcRom[10655] <= 10'b0001000101;
    pxcRom[10656] <= 10'b0000110000;
    pxcRom[10657] <= 10'b0000011101;
    pxcRom[10658] <= 10'b0000010110;
    pxcRom[10659] <= 10'b0000011100;
    pxcRom[10660] <= 10'b0000110000;
    pxcRom[10661] <= 10'b0001010011;
    pxcRom[10662] <= 10'b0010000110;
    pxcRom[10663] <= 10'b0011001001;
    pxcRom[10664] <= 10'b0101000101;
    pxcRom[10665] <= 10'b1000101110;
    pxcRom[10666] <= 10'b1000000001;
    pxcRom[10667] <= 10'b1000101110;
    pxcRom[10668] <= 10'b1000101110;
    pxcRom[10669] <= 10'b0111010101;
    pxcRom[10670] <= 10'b0101000011;
    pxcRom[10671] <= 10'b0011101001;
    pxcRom[10672] <= 10'b0011000010;
    pxcRom[10673] <= 10'b0010101101;
    pxcRom[10674] <= 10'b0010100101;
    pxcRom[10675] <= 10'b0010011100;
    pxcRom[10676] <= 10'b0010010111;
    pxcRom[10677] <= 10'b0010010110;
    pxcRom[10678] <= 10'b0010010011;
    pxcRom[10679] <= 10'b0010010010;
    pxcRom[10680] <= 10'b0010010001;
    pxcRom[10681] <= 10'b0010001011;
    pxcRom[10682] <= 10'b0001111001;
    pxcRom[10683] <= 10'b0001011010;
    pxcRom[10684] <= 10'b0000111011;
    pxcRom[10685] <= 10'b0000100010;
    pxcRom[10686] <= 10'b0000011000;
    pxcRom[10687] <= 10'b0000011011;
    pxcRom[10688] <= 10'b0000101101;
    pxcRom[10689] <= 10'b0001001110;
    pxcRom[10690] <= 10'b0001111010;
    pxcRom[10691] <= 10'b0010111110;
    pxcRom[10692] <= 10'b0100111011;
    pxcRom[10693] <= 10'b1000101110;
    pxcRom[10694] <= 10'b1000101110;
    pxcRom[10695] <= 10'b1000101110;
    pxcRom[10696] <= 10'b1000101110;
    pxcRom[10697] <= 10'b1000000001;
    pxcRom[10698] <= 10'b0100100101;
    pxcRom[10699] <= 10'b0011000101;
    pxcRom[10700] <= 10'b0010011110;
    pxcRom[10701] <= 10'b0010000110;
    pxcRom[10702] <= 10'b0001111011;
    pxcRom[10703] <= 10'b0001110111;
    pxcRom[10704] <= 10'b0001111100;
    pxcRom[10705] <= 10'b0010001000;
    pxcRom[10706] <= 10'b0010010101;
    pxcRom[10707] <= 10'b0010011110;
    pxcRom[10708] <= 10'b0010100100;
    pxcRom[10709] <= 10'b0010011010;
    pxcRom[10710] <= 10'b0001111100;
    pxcRom[10711] <= 10'b0001010101;
    pxcRom[10712] <= 10'b0000110100;
    pxcRom[10713] <= 10'b0000100000;
    pxcRom[10714] <= 10'b0000010111;
    pxcRom[10715] <= 10'b0000011011;
    pxcRom[10716] <= 10'b0000101110;
    pxcRom[10717] <= 10'b0001001110;
    pxcRom[10718] <= 10'b0001110111;
    pxcRom[10719] <= 10'b0010111110;
    pxcRom[10720] <= 10'b0101000000;
    pxcRom[10721] <= 10'b1000101110;
    pxcRom[10722] <= 10'b1000101110;
    pxcRom[10723] <= 10'b1000101110;
    pxcRom[10724] <= 10'b1000101110;
    pxcRom[10725] <= 10'b0111000111;
    pxcRom[10726] <= 10'b0100001101;
    pxcRom[10727] <= 10'b0010110010;
    pxcRom[10728] <= 10'b0010000011;
    pxcRom[10729] <= 10'b0001101010;
    pxcRom[10730] <= 10'b0001011100;
    pxcRom[10731] <= 10'b0001010110;
    pxcRom[10732] <= 10'b0001010111;
    pxcRom[10733] <= 10'b0001011111;
    pxcRom[10734] <= 10'b0001101011;
    pxcRom[10735] <= 10'b0001111001;
    pxcRom[10736] <= 10'b0001111101;
    pxcRom[10737] <= 10'b0001110000;
    pxcRom[10738] <= 10'b0001010111;
    pxcRom[10739] <= 10'b0000111100;
    pxcRom[10740] <= 10'b0000100110;
    pxcRom[10741] <= 10'b0000011000;
    pxcRom[10742] <= 10'b0000010101;
    pxcRom[10743] <= 10'b0000011101;
    pxcRom[10744] <= 10'b0000110100;
    pxcRom[10745] <= 10'b0001010100;
    pxcRom[10746] <= 10'b0010000001;
    pxcRom[10747] <= 10'b0011001100;
    pxcRom[10748] <= 10'b0101100000;
    pxcRom[10749] <= 10'b1000101110;
    pxcRom[10750] <= 10'b1000101110;
    pxcRom[10751] <= 10'b1000101110;
    pxcRom[10752] <= 10'b1000101110;
    pxcRom[10753] <= 10'b0110111011;
    pxcRom[10754] <= 10'b0100000100;
    pxcRom[10755] <= 10'b0010100110;
    pxcRom[10756] <= 10'b0001111001;
    pxcRom[10757] <= 10'b0001011010;
    pxcRom[10758] <= 10'b0001000111;
    pxcRom[10759] <= 10'b0000111100;
    pxcRom[10760] <= 10'b0000111000;
    pxcRom[10761] <= 10'b0000111001;
    pxcRom[10762] <= 10'b0000111110;
    pxcRom[10763] <= 10'b0001000101;
    pxcRom[10764] <= 10'b0001000101;
    pxcRom[10765] <= 10'b0000111101;
    pxcRom[10766] <= 10'b0000101111;
    pxcRom[10767] <= 10'b0000100001;
    pxcRom[10768] <= 10'b0000010101;
    pxcRom[10769] <= 10'b0000010001;
    pxcRom[10770] <= 10'b0000010110;
    pxcRom[10771] <= 10'b0000100110;
    pxcRom[10772] <= 10'b0000111111;
    pxcRom[10773] <= 10'b0001100011;
    pxcRom[10774] <= 10'b0010010110;
    pxcRom[10775] <= 10'b0011101100;
    pxcRom[10776] <= 10'b0110000101;
    pxcRom[10777] <= 10'b1000101110;
    pxcRom[10778] <= 10'b1000000001;
    pxcRom[10779] <= 10'b1000101110;
    pxcRom[10780] <= 10'b1000101110;
    pxcRom[10781] <= 10'b0110110001;
    pxcRom[10782] <= 10'b0100001010;
    pxcRom[10783] <= 10'b0010101101;
    pxcRom[10784] <= 10'b0001111010;
    pxcRom[10785] <= 10'b0001011000;
    pxcRom[10786] <= 10'b0000111110;
    pxcRom[10787] <= 10'b0000101110;
    pxcRom[10788] <= 10'b0000100011;
    pxcRom[10789] <= 10'b0000011111;
    pxcRom[10790] <= 10'b0000011110;
    pxcRom[10791] <= 10'b0000011110;
    pxcRom[10792] <= 10'b0000011101;
    pxcRom[10793] <= 10'b0000011001;
    pxcRom[10794] <= 10'b0000010011;
    pxcRom[10795] <= 10'b0000001111;
    pxcRom[10796] <= 10'b0000001110;
    pxcRom[10797] <= 10'b0000010011;
    pxcRom[10798] <= 10'b0000100000;
    pxcRom[10799] <= 10'b0000110110;
    pxcRom[10800] <= 10'b0001010100;
    pxcRom[10801] <= 10'b0001111111;
    pxcRom[10802] <= 10'b0010111111;
    pxcRom[10803] <= 10'b0100100011;
    pxcRom[10804] <= 10'b0111000111;
    pxcRom[10805] <= 10'b1000101110;
    pxcRom[10806] <= 10'b1000000001;
    pxcRom[10807] <= 10'b1000101110;
    pxcRom[10808] <= 10'b1000101110;
    pxcRom[10809] <= 10'b1000000001;
    pxcRom[10810] <= 10'b0100011110;
    pxcRom[10811] <= 10'b0011000100;
    pxcRom[10812] <= 10'b0010001100;
    pxcRom[10813] <= 10'b0001100100;
    pxcRom[10814] <= 10'b0001000100;
    pxcRom[10815] <= 10'b0000101101;
    pxcRom[10816] <= 10'b0000011110;
    pxcRom[10817] <= 10'b0000010100;
    pxcRom[10818] <= 10'b0000001111;
    pxcRom[10819] <= 10'b0000001100;
    pxcRom[10820] <= 10'b0000001011;
    pxcRom[10821] <= 10'b0000001010;
    pxcRom[10822] <= 10'b0000001010;
    pxcRom[10823] <= 10'b0000001100;
    pxcRom[10824] <= 10'b0000010011;
    pxcRom[10825] <= 10'b0000100001;
    pxcRom[10826] <= 10'b0000110110;
    pxcRom[10827] <= 10'b0001010100;
    pxcRom[10828] <= 10'b0001111011;
    pxcRom[10829] <= 10'b0010110000;
    pxcRom[10830] <= 10'b0011111010;
    pxcRom[10831] <= 10'b0101101000;
    pxcRom[10832] <= 10'b1000000001;
    pxcRom[10833] <= 10'b1000101110;
    pxcRom[10834] <= 10'b1000101110;
    pxcRom[10835] <= 10'b1000101110;
    pxcRom[10836] <= 10'b1000101110;
    pxcRom[10837] <= 10'b1000101110;
    pxcRom[10838] <= 10'b0101001100;
    pxcRom[10839] <= 10'b0011110010;
    pxcRom[10840] <= 10'b0010101110;
    pxcRom[10841] <= 10'b0010000011;
    pxcRom[10842] <= 10'b0001011110;
    pxcRom[10843] <= 10'b0001000000;
    pxcRom[10844] <= 10'b0000101100;
    pxcRom[10845] <= 10'b0000011101;
    pxcRom[10846] <= 10'b0000010100;
    pxcRom[10847] <= 10'b0000010000;
    pxcRom[10848] <= 10'b0000001110;
    pxcRom[10849] <= 10'b0000001111;
    pxcRom[10850] <= 10'b0000010100;
    pxcRom[10851] <= 10'b0000011101;
    pxcRom[10852] <= 10'b0000101101;
    pxcRom[10853] <= 10'b0001000100;
    pxcRom[10854] <= 10'b0001100010;
    pxcRom[10855] <= 10'b0010000110;
    pxcRom[10856] <= 10'b0010111001;
    pxcRom[10857] <= 10'b0011111101;
    pxcRom[10858] <= 10'b0101010100;
    pxcRom[10859] <= 10'b0111000111;
    pxcRom[10860] <= 10'b1000000001;
    pxcRom[10861] <= 10'b1000101110;
    pxcRom[10862] <= 10'b1000000001;
    pxcRom[10863] <= 10'b1000101110;
    pxcRom[10864] <= 10'b1000101110;
    pxcRom[10865] <= 10'b1000101110;
    pxcRom[10866] <= 10'b0110100001;
    pxcRom[10867] <= 10'b0100110110;
    pxcRom[10868] <= 10'b0011110000;
    pxcRom[10869] <= 10'b0011000000;
    pxcRom[10870] <= 10'b0010011001;
    pxcRom[10871] <= 10'b0001111010;
    pxcRom[10872] <= 10'b0001100001;
    pxcRom[10873] <= 10'b0001010000;
    pxcRom[10874] <= 10'b0001000011;
    pxcRom[10875] <= 10'b0000111100;
    pxcRom[10876] <= 10'b0000111011;
    pxcRom[10877] <= 10'b0000111110;
    pxcRom[10878] <= 10'b0001000111;
    pxcRom[10879] <= 10'b0001010101;
    pxcRom[10880] <= 10'b0001101100;
    pxcRom[10881] <= 10'b0010001010;
    pxcRom[10882] <= 10'b0010101110;
    pxcRom[10883] <= 10'b0011011111;
    pxcRom[10884] <= 10'b0100100000;
    pxcRom[10885] <= 10'b0101101110;
    pxcRom[10886] <= 10'b0110100001;
    pxcRom[10887] <= 10'b0111100111;
    pxcRom[10888] <= 10'b1000101110;
    pxcRom[10889] <= 10'b1000101110;
    pxcRom[10890] <= 10'b1000101110;
    pxcRom[10891] <= 10'b1000101110;
    pxcRom[10892] <= 10'b1000101110;
    pxcRom[10893] <= 10'b1000101110;
    pxcRom[10894] <= 10'b1000000001;
    pxcRom[10895] <= 10'b0111100111;
    pxcRom[10896] <= 10'b0110000000;
    pxcRom[10897] <= 10'b0101010100;
    pxcRom[10898] <= 10'b0100100011;
    pxcRom[10899] <= 10'b0011111101;
    pxcRom[10900] <= 10'b0011100101;
    pxcRom[10901] <= 10'b0011010110;
    pxcRom[10902] <= 10'b0011000101;
    pxcRom[10903] <= 10'b0010111011;
    pxcRom[10904] <= 10'b0010111100;
    pxcRom[10905] <= 10'b0010111110;
    pxcRom[10906] <= 10'b0011001000;
    pxcRom[10907] <= 10'b0011011010;
    pxcRom[10908] <= 10'b0011101101;
    pxcRom[10909] <= 10'b0100001010;
    pxcRom[10910] <= 10'b0100101101;
    pxcRom[10911] <= 10'b0101010100;
    pxcRom[10912] <= 10'b0110000101;
    pxcRom[10913] <= 10'b0111000111;
    pxcRom[10914] <= 10'b0111100111;
    pxcRom[10915] <= 10'b1000101110;
    pxcRom[10916] <= 10'b1000101110;
    pxcRom[10917] <= 10'b1000101110;
    pxcRom[10918] <= 10'b1000101110;
    pxcRom[10919] <= 10'b1000101110;
    pxcRom[10920] <= 10'b1000101110;
    pxcRom[10921] <= 10'b1000101110;
    pxcRom[10922] <= 10'b1000101110;
    pxcRom[10923] <= 10'b1000101110;
    pxcRom[10924] <= 10'b1000101110;
    pxcRom[10925] <= 10'b0111100111;
    pxcRom[10926] <= 10'b0111100111;
    pxcRom[10927] <= 10'b0111010101;
    pxcRom[10928] <= 10'b0111000111;
    pxcRom[10929] <= 10'b0111000111;
    pxcRom[10930] <= 10'b0110011010;
    pxcRom[10931] <= 10'b0110010100;
    pxcRom[10932] <= 10'b0110010100;
    pxcRom[10933] <= 10'b0110001111;
    pxcRom[10934] <= 10'b0110010100;
    pxcRom[10935] <= 10'b0110100001;
    pxcRom[10936] <= 10'b0110011010;
    pxcRom[10937] <= 10'b0110100001;
    pxcRom[10938] <= 10'b0110110001;
    pxcRom[10939] <= 10'b0111000111;
    pxcRom[10940] <= 10'b0111010101;
    pxcRom[10941] <= 10'b0111100111;
    pxcRom[10942] <= 10'b1000000001;
    pxcRom[10943] <= 10'b1000101110;
    pxcRom[10944] <= 10'b1000101110;
    pxcRom[10945] <= 10'b1000101110;
    pxcRom[10946] <= 10'b1000101110;
    pxcRom[10947] <= 10'b1000101110;
    pxcRom[10948] <= 10'b1000101110;
    pxcRom[10949] <= 10'b1000101110;
    pxcRom[10950] <= 10'b1000101110;
    pxcRom[10951] <= 10'b1000101110;
    pxcRom[10952] <= 10'b1000101110;
    pxcRom[10953] <= 10'b1000101110;
    pxcRom[10954] <= 10'b1000101110;
    pxcRom[10955] <= 10'b1000101110;
    pxcRom[10956] <= 10'b1000101110;
    pxcRom[10957] <= 10'b1000101110;
    pxcRom[10958] <= 10'b1000101110;
    pxcRom[10959] <= 10'b1000101110;
    pxcRom[10960] <= 10'b1000101110;
    pxcRom[10961] <= 10'b1000101110;
    pxcRom[10962] <= 10'b1000101110;
    pxcRom[10963] <= 10'b1000101110;
    pxcRom[10964] <= 10'b1000101110;
    pxcRom[10965] <= 10'b1000101110;
    pxcRom[10966] <= 10'b1000101110;
    pxcRom[10967] <= 10'b1000101110;
    pxcRom[10968] <= 10'b1000101110;
    pxcRom[10969] <= 10'b1000101110;
    pxcRom[10970] <= 10'b1000101110;
    pxcRom[10971] <= 10'b1000101110;
    pxcRom[10972] <= 10'b1000101110;
    pxcRom[10973] <= 10'b1000101110;
    pxcRom[10974] <= 10'b1000101110;
    pxcRom[10975] <= 10'b1000101110;
    pxcRom[10976] <= 10'b1000101011;
    pxcRom[10977] <= 10'b1000101011;
    pxcRom[10978] <= 10'b1000101011;
    pxcRom[10979] <= 10'b1000101011;
    pxcRom[10980] <= 10'b1000101011;
    pxcRom[10981] <= 10'b1000101011;
    pxcRom[10982] <= 10'b1000101011;
    pxcRom[10983] <= 10'b1000101011;
    pxcRom[10984] <= 10'b1000101011;
    pxcRom[10985] <= 10'b1000101011;
    pxcRom[10986] <= 10'b1000101011;
    pxcRom[10987] <= 10'b1000101011;
    pxcRom[10988] <= 10'b1000101011;
    pxcRom[10989] <= 10'b1000101011;
    pxcRom[10990] <= 10'b1000101011;
    pxcRom[10991] <= 10'b1000101011;
    pxcRom[10992] <= 10'b1000101011;
    pxcRom[10993] <= 10'b1000101011;
    pxcRom[10994] <= 10'b1000101011;
    pxcRom[10995] <= 10'b1000101011;
    pxcRom[10996] <= 10'b1000101011;
    pxcRom[10997] <= 10'b1000101011;
    pxcRom[10998] <= 10'b1000101011;
    pxcRom[10999] <= 10'b1000101011;
    pxcRom[11000] <= 10'b1000101011;
    pxcRom[11001] <= 10'b1000101011;
    pxcRom[11002] <= 10'b1000101011;
    pxcRom[11003] <= 10'b1000101011;
    pxcRom[11004] <= 10'b1000101011;
    pxcRom[11005] <= 10'b1000101011;
    pxcRom[11006] <= 10'b1000101011;
    pxcRom[11007] <= 10'b1000101011;
    pxcRom[11008] <= 10'b1000101011;
    pxcRom[11009] <= 10'b1000101011;
    pxcRom[11010] <= 10'b1000101011;
    pxcRom[11011] <= 10'b1000101011;
    pxcRom[11012] <= 10'b1000101011;
    pxcRom[11013] <= 10'b1000101011;
    pxcRom[11014] <= 10'b1000101011;
    pxcRom[11015] <= 10'b1000101011;
    pxcRom[11016] <= 10'b1000101011;
    pxcRom[11017] <= 10'b1000101011;
    pxcRom[11018] <= 10'b0111111110;
    pxcRom[11019] <= 10'b1000101011;
    pxcRom[11020] <= 10'b1000101011;
    pxcRom[11021] <= 10'b1000101011;
    pxcRom[11022] <= 10'b1000101011;
    pxcRom[11023] <= 10'b1000101011;
    pxcRom[11024] <= 10'b1000101011;
    pxcRom[11025] <= 10'b1000101011;
    pxcRom[11026] <= 10'b1000101011;
    pxcRom[11027] <= 10'b1000101011;
    pxcRom[11028] <= 10'b1000101011;
    pxcRom[11029] <= 10'b1000101011;
    pxcRom[11030] <= 10'b1000101011;
    pxcRom[11031] <= 10'b1000101011;
    pxcRom[11032] <= 10'b1000101011;
    pxcRom[11033] <= 10'b1000101011;
    pxcRom[11034] <= 10'b1000101011;
    pxcRom[11035] <= 10'b1000101011;
    pxcRom[11036] <= 10'b1000101011;
    pxcRom[11037] <= 10'b1000101011;
    pxcRom[11038] <= 10'b1000101011;
    pxcRom[11039] <= 10'b1000101011;
    pxcRom[11040] <= 10'b1000101011;
    pxcRom[11041] <= 10'b1000101011;
    pxcRom[11042] <= 10'b1000101011;
    pxcRom[11043] <= 10'b1000101011;
    pxcRom[11044] <= 10'b0111111110;
    pxcRom[11045] <= 10'b0111010010;
    pxcRom[11046] <= 10'b0111000100;
    pxcRom[11047] <= 10'b0111000100;
    pxcRom[11048] <= 10'b0111010010;
    pxcRom[11049] <= 10'b0111010010;
    pxcRom[11050] <= 10'b1000101011;
    pxcRom[11051] <= 10'b0111100100;
    pxcRom[11052] <= 10'b0111100100;
    pxcRom[11053] <= 10'b0111111110;
    pxcRom[11054] <= 10'b0111111110;
    pxcRom[11055] <= 10'b1000101011;
    pxcRom[11056] <= 10'b1000101011;
    pxcRom[11057] <= 10'b1000101011;
    pxcRom[11058] <= 10'b1000101011;
    pxcRom[11059] <= 10'b1000101011;
    pxcRom[11060] <= 10'b1000101011;
    pxcRom[11061] <= 10'b1000101011;
    pxcRom[11062] <= 10'b1000101011;
    pxcRom[11063] <= 10'b1000101011;
    pxcRom[11064] <= 10'b1000101011;
    pxcRom[11065] <= 10'b1000101011;
    pxcRom[11066] <= 10'b1000101011;
    pxcRom[11067] <= 10'b0111111110;
    pxcRom[11068] <= 10'b0111010010;
    pxcRom[11069] <= 10'b0110100101;
    pxcRom[11070] <= 10'b0110010001;
    pxcRom[11071] <= 10'b0101110101;
    pxcRom[11072] <= 10'b0110000010;
    pxcRom[11073] <= 10'b0101110101;
    pxcRom[11074] <= 10'b0101100101;
    pxcRom[11075] <= 10'b0101010001;
    pxcRom[11076] <= 10'b0101010001;
    pxcRom[11077] <= 10'b0101010001;
    pxcRom[11078] <= 10'b0101001011;
    pxcRom[11079] <= 10'b0100110110;
    pxcRom[11080] <= 10'b0100100101;
    pxcRom[11081] <= 10'b0100101111;
    pxcRom[11082] <= 10'b0101001001;
    pxcRom[11083] <= 10'b0101101110;
    pxcRom[11084] <= 10'b0110011110;
    pxcRom[11085] <= 10'b0111111110;
    pxcRom[11086] <= 10'b1000101011;
    pxcRom[11087] <= 10'b1000101011;
    pxcRom[11088] <= 10'b1000101011;
    pxcRom[11089] <= 10'b1000101011;
    pxcRom[11090] <= 10'b1000101011;
    pxcRom[11091] <= 10'b1000101011;
    pxcRom[11092] <= 10'b0110111000;
    pxcRom[11093] <= 10'b0110000110;
    pxcRom[11094] <= 10'b0101101110;
    pxcRom[11095] <= 10'b0101001011;
    pxcRom[11096] <= 10'b0100101010;
    pxcRom[11097] <= 10'b0100001110;
    pxcRom[11098] <= 10'b0100000010;
    pxcRom[11099] <= 10'b0011110011;
    pxcRom[11100] <= 10'b0011100101;
    pxcRom[11101] <= 10'b0011101010;
    pxcRom[11102] <= 10'b0011110001;
    pxcRom[11103] <= 10'b0011100101;
    pxcRom[11104] <= 10'b0011010010;
    pxcRom[11105] <= 10'b0010111110;
    pxcRom[11106] <= 10'b0010110011;
    pxcRom[11107] <= 10'b0010101001;
    pxcRom[11108] <= 10'b0010100101;
    pxcRom[11109] <= 10'b0010101110;
    pxcRom[11110] <= 10'b0011000100;
    pxcRom[11111] <= 10'b0011100000;
    pxcRom[11112] <= 10'b0100011010;
    pxcRom[11113] <= 10'b0101111001;
    pxcRom[11114] <= 10'b0111111110;
    pxcRom[11115] <= 10'b1000101011;
    pxcRom[11116] <= 10'b1000101011;
    pxcRom[11117] <= 10'b1000101011;
    pxcRom[11118] <= 10'b1000101011;
    pxcRom[11119] <= 10'b0111010010;
    pxcRom[11120] <= 10'b0101100101;
    pxcRom[11121] <= 10'b0100100111;
    pxcRom[11122] <= 10'b0011111001;
    pxcRom[11123] <= 10'b0011011000;
    pxcRom[11124] <= 10'b0010111011;
    pxcRom[11125] <= 10'b0010011111;
    pxcRom[11126] <= 10'b0010010000;
    pxcRom[11127] <= 10'b0010001001;
    pxcRom[11128] <= 10'b0010001000;
    pxcRom[11129] <= 10'b0010010000;
    pxcRom[11130] <= 10'b0010010111;
    pxcRom[11131] <= 10'b0010010101;
    pxcRom[11132] <= 10'b0010000001;
    pxcRom[11133] <= 10'b0001101100;
    pxcRom[11134] <= 10'b0001100000;
    pxcRom[11135] <= 10'b0001011100;
    pxcRom[11136] <= 10'b0001011111;
    pxcRom[11137] <= 10'b0001101010;
    pxcRom[11138] <= 10'b0001111010;
    pxcRom[11139] <= 10'b0010010100;
    pxcRom[11140] <= 10'b0011000000;
    pxcRom[11141] <= 10'b0100100111;
    pxcRom[11142] <= 10'b0111010010;
    pxcRom[11143] <= 10'b1000101011;
    pxcRom[11144] <= 10'b1000101011;
    pxcRom[11145] <= 10'b1000101011;
    pxcRom[11146] <= 10'b1000101011;
    pxcRom[11147] <= 10'b0110010111;
    pxcRom[11148] <= 10'b0100110110;
    pxcRom[11149] <= 10'b0011111011;
    pxcRom[11150] <= 10'b0011001001;
    pxcRom[11151] <= 10'b0010100110;
    pxcRom[11152] <= 10'b0010001000;
    pxcRom[11153] <= 10'b0001101110;
    pxcRom[11154] <= 10'b0001011101;
    pxcRom[11155] <= 10'b0001011000;
    pxcRom[11156] <= 10'b0001011010;
    pxcRom[11157] <= 10'b0001100101;
    pxcRom[11158] <= 10'b0001110011;
    pxcRom[11159] <= 10'b0001110101;
    pxcRom[11160] <= 10'b0001100011;
    pxcRom[11161] <= 10'b0001001101;
    pxcRom[11162] <= 10'b0001000000;
    pxcRom[11163] <= 10'b0000111101;
    pxcRom[11164] <= 10'b0001000010;
    pxcRom[11165] <= 10'b0001001111;
    pxcRom[11166] <= 10'b0001100010;
    pxcRom[11167] <= 10'b0001111101;
    pxcRom[11168] <= 10'b0010101011;
    pxcRom[11169] <= 10'b0100001010;
    pxcRom[11170] <= 10'b0110010111;
    pxcRom[11171] <= 10'b1000101011;
    pxcRom[11172] <= 10'b1000101011;
    pxcRom[11173] <= 10'b1000101011;
    pxcRom[11174] <= 10'b1000101011;
    pxcRom[11175] <= 10'b0101110101;
    pxcRom[11176] <= 10'b0100011001;
    pxcRom[11177] <= 10'b0011011110;
    pxcRom[11178] <= 10'b0010110010;
    pxcRom[11179] <= 10'b0010001010;
    pxcRom[11180] <= 10'b0001101000;
    pxcRom[11181] <= 10'b0001010001;
    pxcRom[11182] <= 10'b0001000100;
    pxcRom[11183] <= 10'b0000111111;
    pxcRom[11184] <= 10'b0001000100;
    pxcRom[11185] <= 10'b0001001111;
    pxcRom[11186] <= 10'b0001100010;
    pxcRom[11187] <= 10'b0001101001;
    pxcRom[11188] <= 10'b0001010101;
    pxcRom[11189] <= 10'b0000111110;
    pxcRom[11190] <= 10'b0000101111;
    pxcRom[11191] <= 10'b0000101110;
    pxcRom[11192] <= 10'b0000110110;
    pxcRom[11193] <= 10'b0001000110;
    pxcRom[11194] <= 10'b0001011110;
    pxcRom[11195] <= 10'b0001111110;
    pxcRom[11196] <= 10'b0010101111;
    pxcRom[11197] <= 10'b0100000110;
    pxcRom[11198] <= 10'b0101111101;
    pxcRom[11199] <= 10'b1000101011;
    pxcRom[11200] <= 10'b1000101011;
    pxcRom[11201] <= 10'b1000101011;
    pxcRom[11202] <= 10'b0111111110;
    pxcRom[11203] <= 10'b0101011111;
    pxcRom[11204] <= 10'b0100000111;
    pxcRom[11205] <= 10'b0011010000;
    pxcRom[11206] <= 10'b0010100000;
    pxcRom[11207] <= 10'b0001110110;
    pxcRom[11208] <= 10'b0001010110;
    pxcRom[11209] <= 10'b0000111110;
    pxcRom[11210] <= 10'b0000110010;
    pxcRom[11211] <= 10'b0000101111;
    pxcRom[11212] <= 10'b0000110101;
    pxcRom[11213] <= 10'b0001000111;
    pxcRom[11214] <= 10'b0001011101;
    pxcRom[11215] <= 10'b0001100100;
    pxcRom[11216] <= 10'b0001001101;
    pxcRom[11217] <= 10'b0000110011;
    pxcRom[11218] <= 10'b0000100100;
    pxcRom[11219] <= 10'b0000100100;
    pxcRom[11220] <= 10'b0000110000;
    pxcRom[11221] <= 10'b0001000110;
    pxcRom[11222] <= 10'b0001100100;
    pxcRom[11223] <= 10'b0010001010;
    pxcRom[11224] <= 10'b0011001001;
    pxcRom[11225] <= 10'b0100100101;
    pxcRom[11226] <= 10'b0110100101;
    pxcRom[11227] <= 10'b1000101011;
    pxcRom[11228] <= 10'b1000101011;
    pxcRom[11229] <= 10'b1000101011;
    pxcRom[11230] <= 10'b0111111110;
    pxcRom[11231] <= 10'b0101100101;
    pxcRom[11232] <= 10'b0100000000;
    pxcRom[11233] <= 10'b0011000110;
    pxcRom[11234] <= 10'b0010010001;
    pxcRom[11235] <= 10'b0001100101;
    pxcRom[11236] <= 10'b0001000110;
    pxcRom[11237] <= 10'b0000101111;
    pxcRom[11238] <= 10'b0000100101;
    pxcRom[11239] <= 10'b0000100101;
    pxcRom[11240] <= 10'b0000110001;
    pxcRom[11241] <= 10'b0001001000;
    pxcRom[11242] <= 10'b0001100101;
    pxcRom[11243] <= 10'b0001100111;
    pxcRom[11244] <= 10'b0001000110;
    pxcRom[11245] <= 10'b0000101000;
    pxcRom[11246] <= 10'b0000011011;
    pxcRom[11247] <= 10'b0000011110;
    pxcRom[11248] <= 10'b0000101111;
    pxcRom[11249] <= 10'b0001001101;
    pxcRom[11250] <= 10'b0001110000;
    pxcRom[11251] <= 10'b0010100111;
    pxcRom[11252] <= 10'b0011110100;
    pxcRom[11253] <= 10'b0101000111;
    pxcRom[11254] <= 10'b0111010010;
    pxcRom[11255] <= 10'b1000101011;
    pxcRom[11256] <= 10'b1000101011;
    pxcRom[11257] <= 10'b1000101011;
    pxcRom[11258] <= 10'b0111100100;
    pxcRom[11259] <= 10'b0101010101;
    pxcRom[11260] <= 10'b0011110011;
    pxcRom[11261] <= 10'b0010110110;
    pxcRom[11262] <= 10'b0010000010;
    pxcRom[11263] <= 10'b0001010111;
    pxcRom[11264] <= 10'b0000110110;
    pxcRom[11265] <= 10'b0000100010;
    pxcRom[11266] <= 10'b0000011100;
    pxcRom[11267] <= 10'b0000100010;
    pxcRom[11268] <= 10'b0000110100;
    pxcRom[11269] <= 10'b0001010011;
    pxcRom[11270] <= 10'b0001111001;
    pxcRom[11271] <= 10'b0001101000;
    pxcRom[11272] <= 10'b0000111011;
    pxcRom[11273] <= 10'b0000011110;
    pxcRom[11274] <= 10'b0000010100;
    pxcRom[11275] <= 10'b0000011100;
    pxcRom[11276] <= 10'b0000110011;
    pxcRom[11277] <= 10'b0001011000;
    pxcRom[11278] <= 10'b0010000110;
    pxcRom[11279] <= 10'b0011001001;
    pxcRom[11280] <= 10'b0100100011;
    pxcRom[11281] <= 10'b0101110101;
    pxcRom[11282] <= 10'b1000101011;
    pxcRom[11283] <= 10'b1000101011;
    pxcRom[11284] <= 10'b1000101011;
    pxcRom[11285] <= 10'b1000101011;
    pxcRom[11286] <= 10'b0111010010;
    pxcRom[11287] <= 10'b0101000111;
    pxcRom[11288] <= 10'b0011101101;
    pxcRom[11289] <= 10'b0010101000;
    pxcRom[11290] <= 10'b0001110000;
    pxcRom[11291] <= 10'b0001000101;
    pxcRom[11292] <= 10'b0000101000;
    pxcRom[11293] <= 10'b0000011000;
    pxcRom[11294] <= 10'b0000010111;
    pxcRom[11295] <= 10'b0000100100;
    pxcRom[11296] <= 10'b0000111111;
    pxcRom[11297] <= 10'b0001101011;
    pxcRom[11298] <= 10'b0010001010;
    pxcRom[11299] <= 10'b0001011110;
    pxcRom[11300] <= 10'b0000101100;
    pxcRom[11301] <= 10'b0000010100;
    pxcRom[11302] <= 10'b0000010000;
    pxcRom[11303] <= 10'b0000011110;
    pxcRom[11304] <= 10'b0000111100;
    pxcRom[11305] <= 10'b0001101000;
    pxcRom[11306] <= 10'b0010011111;
    pxcRom[11307] <= 10'b0011101001;
    pxcRom[11308] <= 10'b0100111110;
    pxcRom[11309] <= 10'b0110011110;
    pxcRom[11310] <= 10'b0111100100;
    pxcRom[11311] <= 10'b1000101011;
    pxcRom[11312] <= 10'b1000101011;
    pxcRom[11313] <= 10'b0111111110;
    pxcRom[11314] <= 10'b0111010010;
    pxcRom[11315] <= 10'b0101000000;
    pxcRom[11316] <= 10'b0011100010;
    pxcRom[11317] <= 10'b0010011001;
    pxcRom[11318] <= 10'b0001011110;
    pxcRom[11319] <= 10'b0000110101;
    pxcRom[11320] <= 10'b0000011100;
    pxcRom[11321] <= 10'b0000010001;
    pxcRom[11322] <= 10'b0000010101;
    pxcRom[11323] <= 10'b0000101000;
    pxcRom[11324] <= 10'b0001001010;
    pxcRom[11325] <= 10'b0001110000;
    pxcRom[11326] <= 10'b0001110011;
    pxcRom[11327] <= 10'b0001000101;
    pxcRom[11328] <= 10'b0000011101;
    pxcRom[11329] <= 10'b0000001101;
    pxcRom[11330] <= 10'b0000001111;
    pxcRom[11331] <= 10'b0000100001;
    pxcRom[11332] <= 10'b0001000011;
    pxcRom[11333] <= 10'b0001110000;
    pxcRom[11334] <= 10'b0010100100;
    pxcRom[11335] <= 10'b0011100011;
    pxcRom[11336] <= 10'b0100011110;
    pxcRom[11337] <= 10'b0101110101;
    pxcRom[11338] <= 10'b0111010010;
    pxcRom[11339] <= 10'b1000101011;
    pxcRom[11340] <= 10'b1000101011;
    pxcRom[11341] <= 10'b0111111110;
    pxcRom[11342] <= 10'b0111100100;
    pxcRom[11343] <= 10'b0100111010;
    pxcRom[11344] <= 10'b0011010010;
    pxcRom[11345] <= 10'b0010000100;
    pxcRom[11346] <= 10'b0001001100;
    pxcRom[11347] <= 10'b0000101000;
    pxcRom[11348] <= 10'b0000010011;
    pxcRom[11349] <= 10'b0000001100;
    pxcRom[11350] <= 10'b0000010011;
    pxcRom[11351] <= 10'b0000100110;
    pxcRom[11352] <= 10'b0000111111;
    pxcRom[11353] <= 10'b0001001110;
    pxcRom[11354] <= 10'b0001000100;
    pxcRom[11355] <= 10'b0000100111;
    pxcRom[11356] <= 10'b0000010000;
    pxcRom[11357] <= 10'b0000001000;
    pxcRom[11358] <= 10'b0000001110;
    pxcRom[11359] <= 10'b0000100010;
    pxcRom[11360] <= 10'b0001000001;
    pxcRom[11361] <= 10'b0001100111;
    pxcRom[11362] <= 10'b0010010100;
    pxcRom[11363] <= 10'b0011000010;
    pxcRom[11364] <= 10'b0011111010;
    pxcRom[11365] <= 10'b0101011010;
    pxcRom[11366] <= 10'b0111000100;
    pxcRom[11367] <= 10'b1000101011;
    pxcRom[11368] <= 10'b1000101011;
    pxcRom[11369] <= 10'b0111111110;
    pxcRom[11370] <= 10'b0111111110;
    pxcRom[11371] <= 10'b0100100110;
    pxcRom[11372] <= 10'b0011000000;
    pxcRom[11373] <= 10'b0001110001;
    pxcRom[11374] <= 10'b0000111110;
    pxcRom[11375] <= 10'b0000011111;
    pxcRom[11376] <= 10'b0000001110;
    pxcRom[11377] <= 10'b0000001001;
    pxcRom[11378] <= 10'b0000001110;
    pxcRom[11379] <= 10'b0000011001;
    pxcRom[11380] <= 10'b0000100010;
    pxcRom[11381] <= 10'b0000100100;
    pxcRom[11382] <= 10'b0000011110;
    pxcRom[11383] <= 10'b0000010001;
    pxcRom[11384] <= 10'b0000000111;
    pxcRom[11385] <= 10'b0000000101;
    pxcRom[11386] <= 10'b0000001101;
    pxcRom[11387] <= 10'b0000011111;
    pxcRom[11388] <= 10'b0000111010;
    pxcRom[11389] <= 10'b0001011011;
    pxcRom[11390] <= 10'b0010000001;
    pxcRom[11391] <= 10'b0010101000;
    pxcRom[11392] <= 10'b0011100001;
    pxcRom[11393] <= 10'b0101001001;
    pxcRom[11394] <= 10'b0111010010;
    pxcRom[11395] <= 10'b1000101011;
    pxcRom[11396] <= 10'b1000101011;
    pxcRom[11397] <= 10'b1000101011;
    pxcRom[11398] <= 10'b0110111000;
    pxcRom[11399] <= 10'b0100011100;
    pxcRom[11400] <= 10'b0010111010;
    pxcRom[11401] <= 10'b0001101000;
    pxcRom[11402] <= 10'b0000111010;
    pxcRom[11403] <= 10'b0000011110;
    pxcRom[11404] <= 10'b0000001111;
    pxcRom[11405] <= 10'b0000001010;
    pxcRom[11406] <= 10'b0000001010;
    pxcRom[11407] <= 10'b0000001110;
    pxcRom[11408] <= 10'b0000001111;
    pxcRom[11409] <= 10'b0000001111;
    pxcRom[11410] <= 10'b0000001100;
    pxcRom[11411] <= 10'b0000000111;
    pxcRom[11412] <= 10'b0000000100;
    pxcRom[11413] <= 10'b0000000100;
    pxcRom[11414] <= 10'b0000001101;
    pxcRom[11415] <= 10'b0000011111;
    pxcRom[11416] <= 10'b0000111011;
    pxcRom[11417] <= 10'b0001011010;
    pxcRom[11418] <= 10'b0001111101;
    pxcRom[11419] <= 10'b0010100010;
    pxcRom[11420] <= 10'b0011011100;
    pxcRom[11421] <= 10'b0100111011;
    pxcRom[11422] <= 10'b0111000100;
    pxcRom[11423] <= 10'b1000101011;
    pxcRom[11424] <= 10'b1000101011;
    pxcRom[11425] <= 10'b1000101011;
    pxcRom[11426] <= 10'b0111111110;
    pxcRom[11427] <= 10'b0100101110;
    pxcRom[11428] <= 10'b0010111111;
    pxcRom[11429] <= 10'b0001101100;
    pxcRom[11430] <= 10'b0001000010;
    pxcRom[11431] <= 10'b0000101000;
    pxcRom[11432] <= 10'b0000011010;
    pxcRom[11433] <= 10'b0000010011;
    pxcRom[11434] <= 10'b0000010001;
    pxcRom[11435] <= 10'b0000010001;
    pxcRom[11436] <= 10'b0000010000;
    pxcRom[11437] <= 10'b0000001111;
    pxcRom[11438] <= 10'b0000001011;
    pxcRom[11439] <= 10'b0000000111;
    pxcRom[11440] <= 10'b0000000100;
    pxcRom[11441] <= 10'b0000001000;
    pxcRom[11442] <= 10'b0000010101;
    pxcRom[11443] <= 10'b0000101011;
    pxcRom[11444] <= 10'b0001001000;
    pxcRom[11445] <= 10'b0001101000;
    pxcRom[11446] <= 10'b0010001101;
    pxcRom[11447] <= 10'b0010110110;
    pxcRom[11448] <= 10'b0011101011;
    pxcRom[11449] <= 10'b0101001111;
    pxcRom[11450] <= 10'b0111000100;
    pxcRom[11451] <= 10'b1000101011;
    pxcRom[11452] <= 10'b1000101011;
    pxcRom[11453] <= 10'b1000101011;
    pxcRom[11454] <= 10'b0111100100;
    pxcRom[11455] <= 10'b0101001001;
    pxcRom[11456] <= 10'b0011010011;
    pxcRom[11457] <= 10'b0010000010;
    pxcRom[11458] <= 10'b0001011001;
    pxcRom[11459] <= 10'b0001000010;
    pxcRom[11460] <= 10'b0000110100;
    pxcRom[11461] <= 10'b0000101101;
    pxcRom[11462] <= 10'b0000101010;
    pxcRom[11463] <= 10'b0000100111;
    pxcRom[11464] <= 10'b0000100100;
    pxcRom[11465] <= 10'b0000011101;
    pxcRom[11466] <= 10'b0000010100;
    pxcRom[11467] <= 10'b0000001100;
    pxcRom[11468] <= 10'b0000001011;
    pxcRom[11469] <= 10'b0000010011;
    pxcRom[11470] <= 10'b0000100101;
    pxcRom[11471] <= 10'b0001000001;
    pxcRom[11472] <= 10'b0001100010;
    pxcRom[11473] <= 10'b0010000100;
    pxcRom[11474] <= 10'b0010101101;
    pxcRom[11475] <= 10'b0011010111;
    pxcRom[11476] <= 10'b0100010000;
    pxcRom[11477] <= 10'b0101111001;
    pxcRom[11478] <= 10'b0111010010;
    pxcRom[11479] <= 10'b1000101011;
    pxcRom[11480] <= 10'b1000101011;
    pxcRom[11481] <= 10'b1000101011;
    pxcRom[11482] <= 10'b0111000100;
    pxcRom[11483] <= 10'b0101101000;
    pxcRom[11484] <= 10'b0011111100;
    pxcRom[11485] <= 10'b0010101011;
    pxcRom[11486] <= 10'b0010000011;
    pxcRom[11487] <= 10'b0001101101;
    pxcRom[11488] <= 10'b0001100010;
    pxcRom[11489] <= 10'b0001011011;
    pxcRom[11490] <= 10'b0001011000;
    pxcRom[11491] <= 10'b0001010000;
    pxcRom[11492] <= 10'b0001000010;
    pxcRom[11493] <= 10'b0000101111;
    pxcRom[11494] <= 10'b0000011111;
    pxcRom[11495] <= 10'b0000010110;
    pxcRom[11496] <= 10'b0000010110;
    pxcRom[11497] <= 10'b0000100010;
    pxcRom[11498] <= 10'b0000111001;
    pxcRom[11499] <= 10'b0001011010;
    pxcRom[11500] <= 10'b0010000001;
    pxcRom[11501] <= 10'b0010101001;
    pxcRom[11502] <= 10'b0011011011;
    pxcRom[11503] <= 10'b0100001001;
    pxcRom[11504] <= 10'b0101010001;
    pxcRom[11505] <= 10'b0110011110;
    pxcRom[11506] <= 10'b0111111110;
    pxcRom[11507] <= 10'b1000101011;
    pxcRom[11508] <= 10'b1000101011;
    pxcRom[11509] <= 10'b1000101011;
    pxcRom[11510] <= 10'b0111111110;
    pxcRom[11511] <= 10'b0110000010;
    pxcRom[11512] <= 10'b0100110000;
    pxcRom[11513] <= 10'b0011100111;
    pxcRom[11514] <= 10'b0011000001;
    pxcRom[11515] <= 10'b0010101101;
    pxcRom[11516] <= 10'b0010100010;
    pxcRom[11517] <= 10'b0010011010;
    pxcRom[11518] <= 10'b0010001001;
    pxcRom[11519] <= 10'b0001110000;
    pxcRom[11520] <= 10'b0001010010;
    pxcRom[11521] <= 10'b0000111000;
    pxcRom[11522] <= 10'b0000100110;
    pxcRom[11523] <= 10'b0000011111;
    pxcRom[11524] <= 10'b0000100001;
    pxcRom[11525] <= 10'b0000101111;
    pxcRom[11526] <= 10'b0001001000;
    pxcRom[11527] <= 10'b0001101001;
    pxcRom[11528] <= 10'b0010010000;
    pxcRom[11529] <= 10'b0010111101;
    pxcRom[11530] <= 10'b0011110001;
    pxcRom[11531] <= 10'b0100101111;
    pxcRom[11532] <= 10'b0110001100;
    pxcRom[11533] <= 10'b0111010010;
    pxcRom[11534] <= 10'b1000101011;
    pxcRom[11535] <= 10'b1000101011;
    pxcRom[11536] <= 10'b1000101011;
    pxcRom[11537] <= 10'b1000101011;
    pxcRom[11538] <= 10'b0111111110;
    pxcRom[11539] <= 10'b0110111000;
    pxcRom[11540] <= 10'b0101100101;
    pxcRom[11541] <= 10'b0100100011;
    pxcRom[11542] <= 10'b0100001000;
    pxcRom[11543] <= 10'b0011111010;
    pxcRom[11544] <= 10'b0011100000;
    pxcRom[11545] <= 10'b0011000000;
    pxcRom[11546] <= 10'b0010011010;
    pxcRom[11547] <= 10'b0001110000;
    pxcRom[11548] <= 10'b0001010000;
    pxcRom[11549] <= 10'b0000111001;
    pxcRom[11550] <= 10'b0000101100;
    pxcRom[11551] <= 10'b0000100111;
    pxcRom[11552] <= 10'b0000101011;
    pxcRom[11553] <= 10'b0000111000;
    pxcRom[11554] <= 10'b0001001111;
    pxcRom[11555] <= 10'b0001101111;
    pxcRom[11556] <= 10'b0010010101;
    pxcRom[11557] <= 10'b0011000001;
    pxcRom[11558] <= 10'b0011110010;
    pxcRom[11559] <= 10'b0100101110;
    pxcRom[11560] <= 10'b0101110101;
    pxcRom[11561] <= 10'b0111100100;
    pxcRom[11562] <= 10'b1000101011;
    pxcRom[11563] <= 10'b1000101011;
    pxcRom[11564] <= 10'b1000101011;
    pxcRom[11565] <= 10'b1000101011;
    pxcRom[11566] <= 10'b1000101011;
    pxcRom[11567] <= 10'b0111100100;
    pxcRom[11568] <= 10'b0110111000;
    pxcRom[11569] <= 10'b0101111001;
    pxcRom[11570] <= 10'b0101010001;
    pxcRom[11571] <= 10'b0100011011;
    pxcRom[11572] <= 10'b0011100001;
    pxcRom[11573] <= 10'b0010110101;
    pxcRom[11574] <= 10'b0010000111;
    pxcRom[11575] <= 10'b0001100101;
    pxcRom[11576] <= 10'b0001001010;
    pxcRom[11577] <= 10'b0000111010;
    pxcRom[11578] <= 10'b0000110010;
    pxcRom[11579] <= 10'b0000101110;
    pxcRom[11580] <= 10'b0000110011;
    pxcRom[11581] <= 10'b0000111111;
    pxcRom[11582] <= 10'b0001010011;
    pxcRom[11583] <= 10'b0001101111;
    pxcRom[11584] <= 10'b0010010010;
    pxcRom[11585] <= 10'b0010111010;
    pxcRom[11586] <= 10'b0011101011;
    pxcRom[11587] <= 10'b0100100001;
    pxcRom[11588] <= 10'b0101100101;
    pxcRom[11589] <= 10'b0111010010;
    pxcRom[11590] <= 10'b1000101011;
    pxcRom[11591] <= 10'b1000101011;
    pxcRom[11592] <= 10'b1000101011;
    pxcRom[11593] <= 10'b1000101011;
    pxcRom[11594] <= 10'b1000101011;
    pxcRom[11595] <= 10'b1000101011;
    pxcRom[11596] <= 10'b1000101011;
    pxcRom[11597] <= 10'b0110011110;
    pxcRom[11598] <= 10'b0101010011;
    pxcRom[11599] <= 10'b0100001101;
    pxcRom[11600] <= 10'b0011010011;
    pxcRom[11601] <= 10'b0010100011;
    pxcRom[11602] <= 10'b0001111011;
    pxcRom[11603] <= 10'b0001011101;
    pxcRom[11604] <= 10'b0001001000;
    pxcRom[11605] <= 10'b0000111110;
    pxcRom[11606] <= 10'b0000111000;
    pxcRom[11607] <= 10'b0000110110;
    pxcRom[11608] <= 10'b0000111001;
    pxcRom[11609] <= 10'b0001000100;
    pxcRom[11610] <= 10'b0001010111;
    pxcRom[11611] <= 10'b0001110000;
    pxcRom[11612] <= 10'b0010010000;
    pxcRom[11613] <= 10'b0010110111;
    pxcRom[11614] <= 10'b0011100100;
    pxcRom[11615] <= 10'b0100011101;
    pxcRom[11616] <= 10'b0101100101;
    pxcRom[11617] <= 10'b0111000100;
    pxcRom[11618] <= 10'b0111111110;
    pxcRom[11619] <= 10'b1000101011;
    pxcRom[11620] <= 10'b1000101011;
    pxcRom[11621] <= 10'b1000101011;
    pxcRom[11622] <= 10'b1000101011;
    pxcRom[11623] <= 10'b1000101011;
    pxcRom[11624] <= 10'b1000101011;
    pxcRom[11625] <= 10'b0111010010;
    pxcRom[11626] <= 10'b0101001001;
    pxcRom[11627] <= 10'b0100000001;
    pxcRom[11628] <= 10'b0011001001;
    pxcRom[11629] <= 10'b0010011100;
    pxcRom[11630] <= 10'b0001111000;
    pxcRom[11631] <= 10'b0001011111;
    pxcRom[11632] <= 10'b0001001111;
    pxcRom[11633] <= 10'b0001000110;
    pxcRom[11634] <= 10'b0001000010;
    pxcRom[11635] <= 10'b0000111111;
    pxcRom[11636] <= 10'b0001000011;
    pxcRom[11637] <= 10'b0001001100;
    pxcRom[11638] <= 10'b0001011101;
    pxcRom[11639] <= 10'b0001110100;
    pxcRom[11640] <= 10'b0010010010;
    pxcRom[11641] <= 10'b0010111100;
    pxcRom[11642] <= 10'b0011101110;
    pxcRom[11643] <= 10'b0100101000;
    pxcRom[11644] <= 10'b0101110010;
    pxcRom[11645] <= 10'b0111010010;
    pxcRom[11646] <= 10'b0111111110;
    pxcRom[11647] <= 10'b1000101011;
    pxcRom[11648] <= 10'b1000101011;
    pxcRom[11649] <= 10'b1000101011;
    pxcRom[11650] <= 10'b1000101011;
    pxcRom[11651] <= 10'b1000101011;
    pxcRom[11652] <= 10'b1000101011;
    pxcRom[11653] <= 10'b0110101110;
    pxcRom[11654] <= 10'b0101001011;
    pxcRom[11655] <= 10'b0100001000;
    pxcRom[11656] <= 10'b0011010111;
    pxcRom[11657] <= 10'b0010101011;
    pxcRom[11658] <= 10'b0010001101;
    pxcRom[11659] <= 10'b0001110101;
    pxcRom[11660] <= 10'b0001100111;
    pxcRom[11661] <= 10'b0001011111;
    pxcRom[11662] <= 10'b0001011011;
    pxcRom[11663] <= 10'b0001011000;
    pxcRom[11664] <= 10'b0001011100;
    pxcRom[11665] <= 10'b0001100111;
    pxcRom[11666] <= 10'b0001110110;
    pxcRom[11667] <= 10'b0010001111;
    pxcRom[11668] <= 10'b0010101011;
    pxcRom[11669] <= 10'b0011011001;
    pxcRom[11670] <= 10'b0100001010;
    pxcRom[11671] <= 10'b0101000011;
    pxcRom[11672] <= 10'b0110100101;
    pxcRom[11673] <= 10'b0111100100;
    pxcRom[11674] <= 10'b1000101011;
    pxcRom[11675] <= 10'b1000101011;
    pxcRom[11676] <= 10'b1000101011;
    pxcRom[11677] <= 10'b1000101011;
    pxcRom[11678] <= 10'b1000101011;
    pxcRom[11679] <= 10'b1000101011;
    pxcRom[11680] <= 10'b0111111110;
    pxcRom[11681] <= 10'b0111100100;
    pxcRom[11682] <= 10'b0110010111;
    pxcRom[11683] <= 10'b0101010001;
    pxcRom[11684] <= 10'b0100011101;
    pxcRom[11685] <= 10'b0011110001;
    pxcRom[11686] <= 10'b0011010111;
    pxcRom[11687] <= 10'b0011000111;
    pxcRom[11688] <= 10'b0010111110;
    pxcRom[11689] <= 10'b0010110000;
    pxcRom[11690] <= 10'b0010100110;
    pxcRom[11691] <= 10'b0010100110;
    pxcRom[11692] <= 10'b0010110000;
    pxcRom[11693] <= 10'b0011000010;
    pxcRom[11694] <= 10'b0011011000;
    pxcRom[11695] <= 10'b0011111001;
    pxcRom[11696] <= 10'b0100011110;
    pxcRom[11697] <= 10'b0101001001;
    pxcRom[11698] <= 10'b0101110010;
    pxcRom[11699] <= 10'b0110001100;
    pxcRom[11700] <= 10'b0111100100;
    pxcRom[11701] <= 10'b1000101011;
    pxcRom[11702] <= 10'b1000101011;
    pxcRom[11703] <= 10'b1000101011;
    pxcRom[11704] <= 10'b1000101011;
    pxcRom[11705] <= 10'b1000101011;
    pxcRom[11706] <= 10'b1000101011;
    pxcRom[11707] <= 10'b1000101011;
    pxcRom[11708] <= 10'b0111111110;
    pxcRom[11709] <= 10'b0111111110;
    pxcRom[11710] <= 10'b0111111110;
    pxcRom[11711] <= 10'b0111111110;
    pxcRom[11712] <= 10'b0111010010;
    pxcRom[11713] <= 10'b0110011110;
    pxcRom[11714] <= 10'b0110001100;
    pxcRom[11715] <= 10'b0101110101;
    pxcRom[11716] <= 10'b0101111001;
    pxcRom[11717] <= 10'b0101101110;
    pxcRom[11718] <= 10'b0101111001;
    pxcRom[11719] <= 10'b0110010001;
    pxcRom[11720] <= 10'b0110010111;
    pxcRom[11721] <= 10'b0110010111;
    pxcRom[11722] <= 10'b0110100101;
    pxcRom[11723] <= 10'b0111010010;
    pxcRom[11724] <= 10'b0111111110;
    pxcRom[11725] <= 10'b1000101011;
    pxcRom[11726] <= 10'b0111111110;
    pxcRom[11727] <= 10'b0111111110;
    pxcRom[11728] <= 10'b1000101011;
    pxcRom[11729] <= 10'b1000101011;
    pxcRom[11730] <= 10'b1000101011;
    pxcRom[11731] <= 10'b1000101011;
    pxcRom[11732] <= 10'b1000101011;
    pxcRom[11733] <= 10'b1000101011;
    pxcRom[11734] <= 10'b1000101011;
    pxcRom[11735] <= 10'b1000101011;
    pxcRom[11736] <= 10'b1000101011;
    pxcRom[11737] <= 10'b1000101011;
    pxcRom[11738] <= 10'b1000101011;
    pxcRom[11739] <= 10'b1000101011;
    pxcRom[11740] <= 10'b1000101011;
    pxcRom[11741] <= 10'b1000101011;
    pxcRom[11742] <= 10'b1000101011;
    pxcRom[11743] <= 10'b1000101011;
    pxcRom[11744] <= 10'b1000101011;
    pxcRom[11745] <= 10'b1000101011;
    pxcRom[11746] <= 10'b1000101011;
    pxcRom[11747] <= 10'b1000101011;
    pxcRom[11748] <= 10'b1000101011;
    pxcRom[11749] <= 10'b1000101011;
    pxcRom[11750] <= 10'b1000101011;
    pxcRom[11751] <= 10'b1000101011;
    pxcRom[11752] <= 10'b1000101011;
    pxcRom[11753] <= 10'b1000101011;
    pxcRom[11754] <= 10'b1000101011;
    pxcRom[11755] <= 10'b1000101011;
    pxcRom[11756] <= 10'b1000101011;
    pxcRom[11757] <= 10'b1000101011;
    pxcRom[11758] <= 10'b1000101011;
    pxcRom[11759] <= 10'b1000101011;
    pxcRom[11760] <= 10'b1000100110;
    pxcRom[11761] <= 10'b1000100110;
    pxcRom[11762] <= 10'b1000100110;
    pxcRom[11763] <= 10'b1000100110;
    pxcRom[11764] <= 10'b1000100110;
    pxcRom[11765] <= 10'b1000100110;
    pxcRom[11766] <= 10'b1000100110;
    pxcRom[11767] <= 10'b1000100110;
    pxcRom[11768] <= 10'b1000100110;
    pxcRom[11769] <= 10'b1000100110;
    pxcRom[11770] <= 10'b1000100110;
    pxcRom[11771] <= 10'b1000100110;
    pxcRom[11772] <= 10'b1000100110;
    pxcRom[11773] <= 10'b1000100110;
    pxcRom[11774] <= 10'b1000100110;
    pxcRom[11775] <= 10'b1000100110;
    pxcRom[11776] <= 10'b1000100110;
    pxcRom[11777] <= 10'b1000100110;
    pxcRom[11778] <= 10'b1000100110;
    pxcRom[11779] <= 10'b1000100110;
    pxcRom[11780] <= 10'b1000100110;
    pxcRom[11781] <= 10'b1000100110;
    pxcRom[11782] <= 10'b1000100110;
    pxcRom[11783] <= 10'b1000100110;
    pxcRom[11784] <= 10'b1000100110;
    pxcRom[11785] <= 10'b1000100110;
    pxcRom[11786] <= 10'b1000100110;
    pxcRom[11787] <= 10'b1000100110;
    pxcRom[11788] <= 10'b1000100110;
    pxcRom[11789] <= 10'b1000100110;
    pxcRom[11790] <= 10'b1000100110;
    pxcRom[11791] <= 10'b1000100110;
    pxcRom[11792] <= 10'b1000100110;
    pxcRom[11793] <= 10'b1000100110;
    pxcRom[11794] <= 10'b1000100110;
    pxcRom[11795] <= 10'b1000100110;
    pxcRom[11796] <= 10'b1000100110;
    pxcRom[11797] <= 10'b1000100110;
    pxcRom[11798] <= 10'b1000100110;
    pxcRom[11799] <= 10'b1000100110;
    pxcRom[11800] <= 10'b1000100110;
    pxcRom[11801] <= 10'b1000100110;
    pxcRom[11802] <= 10'b1000100110;
    pxcRom[11803] <= 10'b1000100110;
    pxcRom[11804] <= 10'b1000100110;
    pxcRom[11805] <= 10'b1000100110;
    pxcRom[11806] <= 10'b1000100110;
    pxcRom[11807] <= 10'b1000100110;
    pxcRom[11808] <= 10'b1000100110;
    pxcRom[11809] <= 10'b1000100110;
    pxcRom[11810] <= 10'b1000100110;
    pxcRom[11811] <= 10'b1000100110;
    pxcRom[11812] <= 10'b1000100110;
    pxcRom[11813] <= 10'b1000100110;
    pxcRom[11814] <= 10'b1000100110;
    pxcRom[11815] <= 10'b1000100110;
    pxcRom[11816] <= 10'b1000100110;
    pxcRom[11817] <= 10'b1000100110;
    pxcRom[11818] <= 10'b1000100110;
    pxcRom[11819] <= 10'b1000100110;
    pxcRom[11820] <= 10'b1000100110;
    pxcRom[11821] <= 10'b1000100110;
    pxcRom[11822] <= 10'b1000100110;
    pxcRom[11823] <= 10'b1000100110;
    pxcRom[11824] <= 10'b1000100110;
    pxcRom[11825] <= 10'b1000100110;
    pxcRom[11826] <= 10'b1000100110;
    pxcRom[11827] <= 10'b1000100110;
    pxcRom[11828] <= 10'b1000100110;
    pxcRom[11829] <= 10'b1000100110;
    pxcRom[11830] <= 10'b0111111001;
    pxcRom[11831] <= 10'b0111001101;
    pxcRom[11832] <= 10'b0110110011;
    pxcRom[11833] <= 10'b0110100001;
    pxcRom[11834] <= 10'b0110100001;
    pxcRom[11835] <= 10'b0110100001;
    pxcRom[11836] <= 10'b0110111111;
    pxcRom[11837] <= 10'b0111011111;
    pxcRom[11838] <= 10'b0111011111;
    pxcRom[11839] <= 10'b0111111001;
    pxcRom[11840] <= 10'b1000100110;
    pxcRom[11841] <= 10'b1000100110;
    pxcRom[11842] <= 10'b1000100110;
    pxcRom[11843] <= 10'b1000100110;
    pxcRom[11844] <= 10'b1000100110;
    pxcRom[11845] <= 10'b1000100110;
    pxcRom[11846] <= 10'b1000100110;
    pxcRom[11847] <= 10'b1000100110;
    pxcRom[11848] <= 10'b0111111001;
    pxcRom[11849] <= 10'b1000100110;
    pxcRom[11850] <= 10'b1000100110;
    pxcRom[11851] <= 10'b1000100110;
    pxcRom[11852] <= 10'b0111111001;
    pxcRom[11853] <= 10'b0110111111;
    pxcRom[11854] <= 10'b0110000111;
    pxcRom[11855] <= 10'b0101101001;
    pxcRom[11856] <= 10'b0101001000;
    pxcRom[11857] <= 10'b0100101110;
    pxcRom[11858] <= 10'b0100011010;
    pxcRom[11859] <= 10'b0100000100;
    pxcRom[11860] <= 10'b0100000110;
    pxcRom[11861] <= 10'b0100000100;
    pxcRom[11862] <= 10'b0100000010;
    pxcRom[11863] <= 10'b0100000100;
    pxcRom[11864] <= 10'b0100001101;
    pxcRom[11865] <= 10'b0100011011;
    pxcRom[11866] <= 10'b0100101001;
    pxcRom[11867] <= 10'b0101011000;
    pxcRom[11868] <= 10'b0101111101;
    pxcRom[11869] <= 10'b0111011111;
    pxcRom[11870] <= 10'b0111111001;
    pxcRom[11871] <= 10'b1000100110;
    pxcRom[11872] <= 10'b1000100110;
    pxcRom[11873] <= 10'b1000100110;
    pxcRom[11874] <= 10'b1000100110;
    pxcRom[11875] <= 10'b1000100110;
    pxcRom[11876] <= 10'b1000100110;
    pxcRom[11877] <= 10'b0111011111;
    pxcRom[11878] <= 10'b0110000010;
    pxcRom[11879] <= 10'b0101001100;
    pxcRom[11880] <= 10'b0100100101;
    pxcRom[11881] <= 10'b0011110001;
    pxcRom[11882] <= 10'b0011001010;
    pxcRom[11883] <= 10'b0010110001;
    pxcRom[11884] <= 10'b0010011111;
    pxcRom[11885] <= 10'b0010001111;
    pxcRom[11886] <= 10'b0010000011;
    pxcRom[11887] <= 10'b0001111100;
    pxcRom[11888] <= 10'b0001110101;
    pxcRom[11889] <= 10'b0001110011;
    pxcRom[11890] <= 10'b0001111000;
    pxcRom[11891] <= 10'b0001111101;
    pxcRom[11892] <= 10'b0010000101;
    pxcRom[11893] <= 10'b0010001101;
    pxcRom[11894] <= 10'b0010011100;
    pxcRom[11895] <= 10'b0010110000;
    pxcRom[11896] <= 10'b0011011000;
    pxcRom[11897] <= 10'b0100011101;
    pxcRom[11898] <= 10'b0110011001;
    pxcRom[11899] <= 10'b1000100110;
    pxcRom[11900] <= 10'b1000100110;
    pxcRom[11901] <= 10'b1000100110;
    pxcRom[11902] <= 10'b1000100110;
    pxcRom[11903] <= 10'b0111111001;
    pxcRom[11904] <= 10'b0111011111;
    pxcRom[11905] <= 10'b0101110000;
    pxcRom[11906] <= 10'b0100011100;
    pxcRom[11907] <= 10'b0011101011;
    pxcRom[11908] <= 10'b0010111111;
    pxcRom[11909] <= 10'b0010011001;
    pxcRom[11910] <= 10'b0001111001;
    pxcRom[11911] <= 10'b0001100001;
    pxcRom[11912] <= 10'b0001010001;
    pxcRom[11913] <= 10'b0001000100;
    pxcRom[11914] <= 10'b0000111101;
    pxcRom[11915] <= 10'b0000111000;
    pxcRom[11916] <= 10'b0000110101;
    pxcRom[11917] <= 10'b0000110101;
    pxcRom[11918] <= 10'b0000110110;
    pxcRom[11919] <= 10'b0000111010;
    pxcRom[11920] <= 10'b0001000000;
    pxcRom[11921] <= 10'b0001001010;
    pxcRom[11922] <= 10'b0001010110;
    pxcRom[11923] <= 10'b0001101001;
    pxcRom[11924] <= 10'b0010000111;
    pxcRom[11925] <= 10'b0011000011;
    pxcRom[11926] <= 10'b0100101001;
    pxcRom[11927] <= 10'b0111011111;
    pxcRom[11928] <= 10'b1000100110;
    pxcRom[11929] <= 10'b1000100110;
    pxcRom[11930] <= 10'b0111111001;
    pxcRom[11931] <= 10'b1000100110;
    pxcRom[11932] <= 10'b0110101001;
    pxcRom[11933] <= 10'b0100101110;
    pxcRom[11934] <= 10'b0011101101;
    pxcRom[11935] <= 10'b0010111100;
    pxcRom[11936] <= 10'b0010010010;
    pxcRom[11937] <= 10'b0001101101;
    pxcRom[11938] <= 10'b0001010011;
    pxcRom[11939] <= 10'b0000111110;
    pxcRom[11940] <= 10'b0000101111;
    pxcRom[11941] <= 10'b0000100110;
    pxcRom[11942] <= 10'b0000100001;
    pxcRom[11943] <= 10'b0000011110;
    pxcRom[11944] <= 10'b0000011110;
    pxcRom[11945] <= 10'b0000011110;
    pxcRom[11946] <= 10'b0000100000;
    pxcRom[11947] <= 10'b0000100100;
    pxcRom[11948] <= 10'b0000101010;
    pxcRom[11949] <= 10'b0000110010;
    pxcRom[11950] <= 10'b0000111100;
    pxcRom[11951] <= 10'b0001001010;
    pxcRom[11952] <= 10'b0001100010;
    pxcRom[11953] <= 10'b0010010101;
    pxcRom[11954] <= 10'b0011110110;
    pxcRom[11955] <= 10'b0110000010;
    pxcRom[11956] <= 10'b1000100110;
    pxcRom[11957] <= 10'b1000100110;
    pxcRom[11958] <= 10'b0111111001;
    pxcRom[11959] <= 10'b1000100110;
    pxcRom[11960] <= 10'b0110101001;
    pxcRom[11961] <= 10'b0100010111;
    pxcRom[11962] <= 10'b0011010001;
    pxcRom[11963] <= 10'b0010011111;
    pxcRom[11964] <= 10'b0001110110;
    pxcRom[11965] <= 10'b0001010101;
    pxcRom[11966] <= 10'b0000111100;
    pxcRom[11967] <= 10'b0000101011;
    pxcRom[11968] <= 10'b0000100000;
    pxcRom[11969] <= 10'b0000011011;
    pxcRom[11970] <= 10'b0000011000;
    pxcRom[11971] <= 10'b0000011000;
    pxcRom[11972] <= 10'b0000011001;
    pxcRom[11973] <= 10'b0000011010;
    pxcRom[11974] <= 10'b0000011101;
    pxcRom[11975] <= 10'b0000100000;
    pxcRom[11976] <= 10'b0000100110;
    pxcRom[11977] <= 10'b0000101101;
    pxcRom[11978] <= 10'b0000110110;
    pxcRom[11979] <= 10'b0001000001;
    pxcRom[11980] <= 10'b0001010101;
    pxcRom[11981] <= 10'b0010000001;
    pxcRom[11982] <= 10'b0011011111;
    pxcRom[11983] <= 10'b0110001100;
    pxcRom[11984] <= 10'b1000100110;
    pxcRom[11985] <= 10'b1000100110;
    pxcRom[11986] <= 10'b1000100110;
    pxcRom[11987] <= 10'b1000100110;
    pxcRom[11988] <= 10'b0110001100;
    pxcRom[11989] <= 10'b0100000100;
    pxcRom[11990] <= 10'b0011000010;
    pxcRom[11991] <= 10'b0010001101;
    pxcRom[11992] <= 10'b0001100011;
    pxcRom[11993] <= 10'b0001000100;
    pxcRom[11994] <= 10'b0000101111;
    pxcRom[11995] <= 10'b0000100000;
    pxcRom[11996] <= 10'b0000011011;
    pxcRom[11997] <= 10'b0000011001;
    pxcRom[11998] <= 10'b0000011011;
    pxcRom[11999] <= 10'b0000011101;
    pxcRom[12000] <= 10'b0000100000;
    pxcRom[12001] <= 10'b0000100011;
    pxcRom[12002] <= 10'b0000101000;
    pxcRom[12003] <= 10'b0000101100;
    pxcRom[12004] <= 10'b0000110010;
    pxcRom[12005] <= 10'b0000111000;
    pxcRom[12006] <= 10'b0001000000;
    pxcRom[12007] <= 10'b0001001010;
    pxcRom[12008] <= 10'b0001011011;
    pxcRom[12009] <= 10'b0010000011;
    pxcRom[12010] <= 10'b0011101000;
    pxcRom[12011] <= 10'b0110100001;
    pxcRom[12012] <= 10'b1000100110;
    pxcRom[12013] <= 10'b1000100110;
    pxcRom[12014] <= 10'b1000100110;
    pxcRom[12015] <= 10'b1000100110;
    pxcRom[12016] <= 10'b0101100110;
    pxcRom[12017] <= 10'b0011110110;
    pxcRom[12018] <= 10'b0010110001;
    pxcRom[12019] <= 10'b0001111100;
    pxcRom[12020] <= 10'b0001010100;
    pxcRom[12021] <= 10'b0000111001;
    pxcRom[12022] <= 10'b0000100101;
    pxcRom[12023] <= 10'b0000011011;
    pxcRom[12024] <= 10'b0000011010;
    pxcRom[12025] <= 10'b0000011110;
    pxcRom[12026] <= 10'b0000100101;
    pxcRom[12027] <= 10'b0000101101;
    pxcRom[12028] <= 10'b0000110011;
    pxcRom[12029] <= 10'b0000111001;
    pxcRom[12030] <= 10'b0000111111;
    pxcRom[12031] <= 10'b0001000100;
    pxcRom[12032] <= 10'b0001001011;
    pxcRom[12033] <= 10'b0001010010;
    pxcRom[12034] <= 10'b0001011010;
    pxcRom[12035] <= 10'b0001100100;
    pxcRom[12036] <= 10'b0001110011;
    pxcRom[12037] <= 10'b0010011010;
    pxcRom[12038] <= 10'b0100000000;
    pxcRom[12039] <= 10'b0110100001;
    pxcRom[12040] <= 10'b1000100110;
    pxcRom[12041] <= 10'b1000100110;
    pxcRom[12042] <= 10'b1000100110;
    pxcRom[12043] <= 10'b1000100110;
    pxcRom[12044] <= 10'b0101000100;
    pxcRom[12045] <= 10'b0011101100;
    pxcRom[12046] <= 10'b0010100011;
    pxcRom[12047] <= 10'b0001101111;
    pxcRom[12048] <= 10'b0001001000;
    pxcRom[12049] <= 10'b0000101100;
    pxcRom[12050] <= 10'b0000011100;
    pxcRom[12051] <= 10'b0000010110;
    pxcRom[12052] <= 10'b0000011001;
    pxcRom[12053] <= 10'b0000100010;
    pxcRom[12054] <= 10'b0000101111;
    pxcRom[12055] <= 10'b0000111011;
    pxcRom[12056] <= 10'b0001001000;
    pxcRom[12057] <= 10'b0001010100;
    pxcRom[12058] <= 10'b0001011111;
    pxcRom[12059] <= 10'b0001101010;
    pxcRom[12060] <= 10'b0001110101;
    pxcRom[12061] <= 10'b0010000000;
    pxcRom[12062] <= 10'b0010001001;
    pxcRom[12063] <= 10'b0010010100;
    pxcRom[12064] <= 10'b0010100011;
    pxcRom[12065] <= 10'b0011001010;
    pxcRom[12066] <= 10'b0100100100;
    pxcRom[12067] <= 10'b0111001101;
    pxcRom[12068] <= 10'b1000100110;
    pxcRom[12069] <= 10'b1000100110;
    pxcRom[12070] <= 10'b1000100110;
    pxcRom[12071] <= 10'b0111001101;
    pxcRom[12072] <= 10'b0100110101;
    pxcRom[12073] <= 10'b0011011101;
    pxcRom[12074] <= 10'b0010011001;
    pxcRom[12075] <= 10'b0001100011;
    pxcRom[12076] <= 10'b0000111101;
    pxcRom[12077] <= 10'b0000100011;
    pxcRom[12078] <= 10'b0000010100;
    pxcRom[12079] <= 10'b0000010001;
    pxcRom[12080] <= 10'b0000010110;
    pxcRom[12081] <= 10'b0000100001;
    pxcRom[12082] <= 10'b0000110000;
    pxcRom[12083] <= 10'b0000111110;
    pxcRom[12084] <= 10'b0001001011;
    pxcRom[12085] <= 10'b0001011100;
    pxcRom[12086] <= 10'b0001101111;
    pxcRom[12087] <= 10'b0010001000;
    pxcRom[12088] <= 10'b0010100001;
    pxcRom[12089] <= 10'b0010111001;
    pxcRom[12090] <= 10'b0011001110;
    pxcRom[12091] <= 10'b0011010111;
    pxcRom[12092] <= 10'b0011100110;
    pxcRom[12093] <= 10'b0100001011;
    pxcRom[12094] <= 10'b0101100000;
    pxcRom[12095] <= 10'b0111111001;
    pxcRom[12096] <= 10'b1000100110;
    pxcRom[12097] <= 10'b1000100110;
    pxcRom[12098] <= 10'b1000100110;
    pxcRom[12099] <= 10'b0110101001;
    pxcRom[12100] <= 10'b0100110001;
    pxcRom[12101] <= 10'b0011010010;
    pxcRom[12102] <= 10'b0010001111;
    pxcRom[12103] <= 10'b0001011010;
    pxcRom[12104] <= 10'b0000110100;
    pxcRom[12105] <= 10'b0000011011;
    pxcRom[12106] <= 10'b0000001110;
    pxcRom[12107] <= 10'b0000001100;
    pxcRom[12108] <= 10'b0000010010;
    pxcRom[12109] <= 10'b0000011100;
    pxcRom[12110] <= 10'b0000100111;
    pxcRom[12111] <= 10'b0000110001;
    pxcRom[12112] <= 10'b0000111101;
    pxcRom[12113] <= 10'b0001001010;
    pxcRom[12114] <= 10'b0001011110;
    pxcRom[12115] <= 10'b0001111100;
    pxcRom[12116] <= 10'b0010011110;
    pxcRom[12117] <= 10'b0011001011;
    pxcRom[12118] <= 10'b0011111010;
    pxcRom[12119] <= 10'b0100011011;
    pxcRom[12120] <= 10'b0101001100;
    pxcRom[12121] <= 10'b0101111000;
    pxcRom[12122] <= 10'b0110110011;
    pxcRom[12123] <= 10'b1000100110;
    pxcRom[12124] <= 10'b1000100110;
    pxcRom[12125] <= 10'b1000100110;
    pxcRom[12126] <= 10'b1000100110;
    pxcRom[12127] <= 10'b0110100001;
    pxcRom[12128] <= 10'b0100101110;
    pxcRom[12129] <= 10'b0011010001;
    pxcRom[12130] <= 10'b0010001110;
    pxcRom[12131] <= 10'b0001011000;
    pxcRom[12132] <= 10'b0000110010;
    pxcRom[12133] <= 10'b0000011001;
    pxcRom[12134] <= 10'b0000001110;
    pxcRom[12135] <= 10'b0000001100;
    pxcRom[12136] <= 10'b0000010000;
    pxcRom[12137] <= 10'b0000010111;
    pxcRom[12138] <= 10'b0000011101;
    pxcRom[12139] <= 10'b0000100100;
    pxcRom[12140] <= 10'b0000101101;
    pxcRom[12141] <= 10'b0000110111;
    pxcRom[12142] <= 10'b0001000101;
    pxcRom[12143] <= 10'b0001011101;
    pxcRom[12144] <= 10'b0001111110;
    pxcRom[12145] <= 10'b0010101101;
    pxcRom[12146] <= 10'b0011100010;
    pxcRom[12147] <= 10'b0100011111;
    pxcRom[12148] <= 10'b0101101101;
    pxcRom[12149] <= 10'b0110111111;
    pxcRom[12150] <= 10'b0111011111;
    pxcRom[12151] <= 10'b1000100110;
    pxcRom[12152] <= 10'b0111111001;
    pxcRom[12153] <= 10'b1000100110;
    pxcRom[12154] <= 10'b1000100110;
    pxcRom[12155] <= 10'b0110101001;
    pxcRom[12156] <= 10'b0100110101;
    pxcRom[12157] <= 10'b0011010111;
    pxcRom[12158] <= 10'b0010010100;
    pxcRom[12159] <= 10'b0001100001;
    pxcRom[12160] <= 10'b0000111010;
    pxcRom[12161] <= 10'b0000100010;
    pxcRom[12162] <= 10'b0000010111;
    pxcRom[12163] <= 10'b0000010101;
    pxcRom[12164] <= 10'b0000010111;
    pxcRom[12165] <= 10'b0000011011;
    pxcRom[12166] <= 10'b0000011110;
    pxcRom[12167] <= 10'b0000100010;
    pxcRom[12168] <= 10'b0000100110;
    pxcRom[12169] <= 10'b0000101100;
    pxcRom[12170] <= 10'b0000110110;
    pxcRom[12171] <= 10'b0001001000;
    pxcRom[12172] <= 10'b0001100100;
    pxcRom[12173] <= 10'b0010001100;
    pxcRom[12174] <= 10'b0010111100;
    pxcRom[12175] <= 10'b0011111101;
    pxcRom[12176] <= 10'b0101010001;
    pxcRom[12177] <= 10'b0111011111;
    pxcRom[12178] <= 10'b1000100110;
    pxcRom[12179] <= 10'b1000100110;
    pxcRom[12180] <= 10'b0111111001;
    pxcRom[12181] <= 10'b1000100110;
    pxcRom[12182] <= 10'b1000100110;
    pxcRom[12183] <= 10'b0110010010;
    pxcRom[12184] <= 10'b0100111010;
    pxcRom[12185] <= 10'b0011011110;
    pxcRom[12186] <= 10'b0010100000;
    pxcRom[12187] <= 10'b0001110011;
    pxcRom[12188] <= 10'b0001001110;
    pxcRom[12189] <= 10'b0000110111;
    pxcRom[12190] <= 10'b0000101101;
    pxcRom[12191] <= 10'b0000101010;
    pxcRom[12192] <= 10'b0000101010;
    pxcRom[12193] <= 10'b0000101011;
    pxcRom[12194] <= 10'b0000101010;
    pxcRom[12195] <= 10'b0000101010;
    pxcRom[12196] <= 10'b0000101000;
    pxcRom[12197] <= 10'b0000101001;
    pxcRom[12198] <= 10'b0000101110;
    pxcRom[12199] <= 10'b0000111100;
    pxcRom[12200] <= 10'b0001010101;
    pxcRom[12201] <= 10'b0001111000;
    pxcRom[12202] <= 10'b0010100010;
    pxcRom[12203] <= 10'b0011010111;
    pxcRom[12204] <= 10'b0100101101;
    pxcRom[12205] <= 10'b0110101001;
    pxcRom[12206] <= 10'b1000100110;
    pxcRom[12207] <= 10'b1000100110;
    pxcRom[12208] <= 10'b1000100110;
    pxcRom[12209] <= 10'b1000100110;
    pxcRom[12210] <= 10'b1000100110;
    pxcRom[12211] <= 10'b0110000010;
    pxcRom[12212] <= 10'b0100011100;
    pxcRom[12213] <= 10'b0011000101;
    pxcRom[12214] <= 10'b0010011011;
    pxcRom[12215] <= 10'b0010000010;
    pxcRom[12216] <= 10'b0001101011;
    pxcRom[12217] <= 10'b0001011001;
    pxcRom[12218] <= 10'b0001010001;
    pxcRom[12219] <= 10'b0001001110;
    pxcRom[12220] <= 10'b0001001011;
    pxcRom[12221] <= 10'b0001000111;
    pxcRom[12222] <= 10'b0000111111;
    pxcRom[12223] <= 10'b0000110110;
    pxcRom[12224] <= 10'b0000101110;
    pxcRom[12225] <= 10'b0000101001;
    pxcRom[12226] <= 10'b0000101011;
    pxcRom[12227] <= 10'b0000110110;
    pxcRom[12228] <= 10'b0001001100;
    pxcRom[12229] <= 10'b0001101011;
    pxcRom[12230] <= 10'b0010010101;
    pxcRom[12231] <= 10'b0011000101;
    pxcRom[12232] <= 10'b0100010010;
    pxcRom[12233] <= 10'b0110110011;
    pxcRom[12234] <= 10'b1000100110;
    pxcRom[12235] <= 10'b1000100110;
    pxcRom[12236] <= 10'b1000100110;
    pxcRom[12237] <= 10'b1000100110;
    pxcRom[12238] <= 10'b1000100110;
    pxcRom[12239] <= 10'b0101110000;
    pxcRom[12240] <= 10'b0011110000;
    pxcRom[12241] <= 10'b0010100000;
    pxcRom[12242] <= 10'b0001111100;
    pxcRom[12243] <= 10'b0001110101;
    pxcRom[12244] <= 10'b0001110110;
    pxcRom[12245] <= 10'b0001110110;
    pxcRom[12246] <= 10'b0001110110;
    pxcRom[12247] <= 10'b0001110101;
    pxcRom[12248] <= 10'b0001110001;
    pxcRom[12249] <= 10'b0001100000;
    pxcRom[12250] <= 10'b0001001110;
    pxcRom[12251] <= 10'b0000111101;
    pxcRom[12252] <= 10'b0000110000;
    pxcRom[12253] <= 10'b0000101001;
    pxcRom[12254] <= 10'b0000101010;
    pxcRom[12255] <= 10'b0000110011;
    pxcRom[12256] <= 10'b0001001000;
    pxcRom[12257] <= 10'b0001100110;
    pxcRom[12258] <= 10'b0010001101;
    pxcRom[12259] <= 10'b0010111100;
    pxcRom[12260] <= 10'b0100000111;
    pxcRom[12261] <= 10'b0110101001;
    pxcRom[12262] <= 10'b0111111001;
    pxcRom[12263] <= 10'b1000100110;
    pxcRom[12264] <= 10'b1000100110;
    pxcRom[12265] <= 10'b1000100110;
    pxcRom[12266] <= 10'b0111111001;
    pxcRom[12267] <= 10'b0101011101;
    pxcRom[12268] <= 10'b0011010000;
    pxcRom[12269] <= 10'b0010000011;
    pxcRom[12270] <= 10'b0001011111;
    pxcRom[12271] <= 10'b0001011010;
    pxcRom[12272] <= 10'b0001100001;
    pxcRom[12273] <= 10'b0001101100;
    pxcRom[12274] <= 10'b0001111010;
    pxcRom[12275] <= 10'b0001111111;
    pxcRom[12276] <= 10'b0001111000;
    pxcRom[12277] <= 10'b0001100101;
    pxcRom[12278] <= 10'b0001001110;
    pxcRom[12279] <= 10'b0000111010;
    pxcRom[12280] <= 10'b0000101101;
    pxcRom[12281] <= 10'b0000100111;
    pxcRom[12282] <= 10'b0000101001;
    pxcRom[12283] <= 10'b0000110100;
    pxcRom[12284] <= 10'b0001001001;
    pxcRom[12285] <= 10'b0001100101;
    pxcRom[12286] <= 10'b0010001010;
    pxcRom[12287] <= 10'b0010111010;
    pxcRom[12288] <= 10'b0100000100;
    pxcRom[12289] <= 10'b0110101001;
    pxcRom[12290] <= 10'b0111111001;
    pxcRom[12291] <= 10'b1000100110;
    pxcRom[12292] <= 10'b1000100110;
    pxcRom[12293] <= 10'b1000100110;
    pxcRom[12294] <= 10'b0111001101;
    pxcRom[12295] <= 10'b0101011010;
    pxcRom[12296] <= 10'b0011000100;
    pxcRom[12297] <= 10'b0001110011;
    pxcRom[12298] <= 10'b0001001100;
    pxcRom[12299] <= 10'b0001000000;
    pxcRom[12300] <= 10'b0001000010;
    pxcRom[12301] <= 10'b0001001100;
    pxcRom[12302] <= 10'b0001010110;
    pxcRom[12303] <= 10'b0001011101;
    pxcRom[12304] <= 10'b0001011010;
    pxcRom[12305] <= 10'b0001001111;
    pxcRom[12306] <= 10'b0000111111;
    pxcRom[12307] <= 10'b0000110000;
    pxcRom[12308] <= 10'b0000100111;
    pxcRom[12309] <= 10'b0000100101;
    pxcRom[12310] <= 10'b0000101000;
    pxcRom[12311] <= 10'b0000110110;
    pxcRom[12312] <= 10'b0001001100;
    pxcRom[12313] <= 10'b0001101001;
    pxcRom[12314] <= 10'b0010001111;
    pxcRom[12315] <= 10'b0011000001;
    pxcRom[12316] <= 10'b0100001111;
    pxcRom[12317] <= 10'b0110011001;
    pxcRom[12318] <= 10'b0111111001;
    pxcRom[12319] <= 10'b1000100110;
    pxcRom[12320] <= 10'b1000100110;
    pxcRom[12321] <= 10'b1000100110;
    pxcRom[12322] <= 10'b0110111111;
    pxcRom[12323] <= 10'b0101001110;
    pxcRom[12324] <= 10'b0011001011;
    pxcRom[12325] <= 10'b0001110100;
    pxcRom[12326] <= 10'b0001000110;
    pxcRom[12327] <= 10'b0000110010;
    pxcRom[12328] <= 10'b0000101100;
    pxcRom[12329] <= 10'b0000101100;
    pxcRom[12330] <= 10'b0000110001;
    pxcRom[12331] <= 10'b0000110110;
    pxcRom[12332] <= 10'b0000110111;
    pxcRom[12333] <= 10'b0000110010;
    pxcRom[12334] <= 10'b0000101010;
    pxcRom[12335] <= 10'b0000100011;
    pxcRom[12336] <= 10'b0000011111;
    pxcRom[12337] <= 10'b0000100001;
    pxcRom[12338] <= 10'b0000101001;
    pxcRom[12339] <= 10'b0000111011;
    pxcRom[12340] <= 10'b0001010011;
    pxcRom[12341] <= 10'b0001110101;
    pxcRom[12342] <= 10'b0010011101;
    pxcRom[12343] <= 10'b0011010101;
    pxcRom[12344] <= 10'b0100100100;
    pxcRom[12345] <= 10'b0110110011;
    pxcRom[12346] <= 10'b0111111001;
    pxcRom[12347] <= 10'b0111111001;
    pxcRom[12348] <= 10'b1000100110;
    pxcRom[12349] <= 10'b1000100110;
    pxcRom[12350] <= 10'b0111111001;
    pxcRom[12351] <= 10'b0101011101;
    pxcRom[12352] <= 10'b0011011110;
    pxcRom[12353] <= 10'b0010000100;
    pxcRom[12354] <= 10'b0001001101;
    pxcRom[12355] <= 10'b0000110001;
    pxcRom[12356] <= 10'b0000100011;
    pxcRom[12357] <= 10'b0000011101;
    pxcRom[12358] <= 10'b0000011100;
    pxcRom[12359] <= 10'b0000011100;
    pxcRom[12360] <= 10'b0000011101;
    pxcRom[12361] <= 10'b0000011100;
    pxcRom[12362] <= 10'b0000011001;
    pxcRom[12363] <= 10'b0000011001;
    pxcRom[12364] <= 10'b0000011011;
    pxcRom[12365] <= 10'b0000100010;
    pxcRom[12366] <= 10'b0000110001;
    pxcRom[12367] <= 10'b0001000111;
    pxcRom[12368] <= 10'b0001100100;
    pxcRom[12369] <= 10'b0010000111;
    pxcRom[12370] <= 10'b0010110110;
    pxcRom[12371] <= 10'b0011110011;
    pxcRom[12372] <= 10'b0101011000;
    pxcRom[12373] <= 10'b0111001101;
    pxcRom[12374] <= 10'b0111111001;
    pxcRom[12375] <= 10'b1000100110;
    pxcRom[12376] <= 10'b1000100110;
    pxcRom[12377] <= 10'b1000100110;
    pxcRom[12378] <= 10'b1000100110;
    pxcRom[12379] <= 10'b0110001100;
    pxcRom[12380] <= 10'b0100000010;
    pxcRom[12381] <= 10'b0010100111;
    pxcRom[12382] <= 10'b0001100111;
    pxcRom[12383] <= 10'b0001000001;
    pxcRom[12384] <= 10'b0000101010;
    pxcRom[12385] <= 10'b0000011100;
    pxcRom[12386] <= 10'b0000010110;
    pxcRom[12387] <= 10'b0000010011;
    pxcRom[12388] <= 10'b0000010010;
    pxcRom[12389] <= 10'b0000010011;
    pxcRom[12390] <= 10'b0000010101;
    pxcRom[12391] <= 10'b0000011000;
    pxcRom[12392] <= 10'b0000100000;
    pxcRom[12393] <= 10'b0000101101;
    pxcRom[12394] <= 10'b0001000001;
    pxcRom[12395] <= 10'b0001011101;
    pxcRom[12396] <= 10'b0001111111;
    pxcRom[12397] <= 10'b0010101011;
    pxcRom[12398] <= 10'b0011011111;
    pxcRom[12399] <= 10'b0100011111;
    pxcRom[12400] <= 10'b0110000010;
    pxcRom[12401] <= 10'b0110111111;
    pxcRom[12402] <= 10'b0111111001;
    pxcRom[12403] <= 10'b1000100110;
    pxcRom[12404] <= 10'b1000100110;
    pxcRom[12405] <= 10'b1000100110;
    pxcRom[12406] <= 10'b0111111001;
    pxcRom[12407] <= 10'b0110100001;
    pxcRom[12408] <= 10'b0100101101;
    pxcRom[12409] <= 10'b0011010111;
    pxcRom[12410] <= 10'b0010010001;
    pxcRom[12411] <= 10'b0001100011;
    pxcRom[12412] <= 10'b0001000100;
    pxcRom[12413] <= 10'b0000110000;
    pxcRom[12414] <= 10'b0000100011;
    pxcRom[12415] <= 10'b0000011100;
    pxcRom[12416] <= 10'b0000011011;
    pxcRom[12417] <= 10'b0000011100;
    pxcRom[12418] <= 10'b0000100000;
    pxcRom[12419] <= 10'b0000101000;
    pxcRom[12420] <= 10'b0000110101;
    pxcRom[12421] <= 10'b0001001010;
    pxcRom[12422] <= 10'b0001100110;
    pxcRom[12423] <= 10'b0010000110;
    pxcRom[12424] <= 10'b0010110010;
    pxcRom[12425] <= 10'b0011100100;
    pxcRom[12426] <= 10'b0100100011;
    pxcRom[12427] <= 10'b0101010011;
    pxcRom[12428] <= 10'b0110110011;
    pxcRom[12429] <= 10'b0111011111;
    pxcRom[12430] <= 10'b0111111001;
    pxcRom[12431] <= 10'b1000100110;
    pxcRom[12432] <= 10'b1000100110;
    pxcRom[12433] <= 10'b1000100110;
    pxcRom[12434] <= 10'b1000100110;
    pxcRom[12435] <= 10'b0111011111;
    pxcRom[12436] <= 10'b0101111101;
    pxcRom[12437] <= 10'b0100101110;
    pxcRom[12438] <= 10'b0011011000;
    pxcRom[12439] <= 10'b0010100010;
    pxcRom[12440] <= 10'b0001111100;
    pxcRom[12441] <= 10'b0001100010;
    pxcRom[12442] <= 10'b0001010000;
    pxcRom[12443] <= 10'b0001000110;
    pxcRom[12444] <= 10'b0001000001;
    pxcRom[12445] <= 10'b0001000011;
    pxcRom[12446] <= 10'b0001001011;
    pxcRom[12447] <= 10'b0001011000;
    pxcRom[12448] <= 10'b0001101101;
    pxcRom[12449] <= 10'b0010001010;
    pxcRom[12450] <= 10'b0010101000;
    pxcRom[12451] <= 10'b0011010001;
    pxcRom[12452] <= 10'b0011111110;
    pxcRom[12453] <= 10'b0100110101;
    pxcRom[12454] <= 10'b0101011101;
    pxcRom[12455] <= 10'b0110011001;
    pxcRom[12456] <= 10'b0111001101;
    pxcRom[12457] <= 10'b1000100110;
    pxcRom[12458] <= 10'b1000100110;
    pxcRom[12459] <= 10'b1000100110;
    pxcRom[12460] <= 10'b1000100110;
    pxcRom[12461] <= 10'b1000100110;
    pxcRom[12462] <= 10'b1000100110;
    pxcRom[12463] <= 10'b0111111001;
    pxcRom[12464] <= 10'b0111011111;
    pxcRom[12465] <= 10'b0110101001;
    pxcRom[12466] <= 10'b0101000110;
    pxcRom[12467] <= 10'b0100010000;
    pxcRom[12468] <= 10'b0011100111;
    pxcRom[12469] <= 10'b0011001010;
    pxcRom[12470] <= 10'b0010111000;
    pxcRom[12471] <= 10'b0010101110;
    pxcRom[12472] <= 10'b0010110000;
    pxcRom[12473] <= 10'b0010110001;
    pxcRom[12474] <= 10'b0011000000;
    pxcRom[12475] <= 10'b0011010001;
    pxcRom[12476] <= 10'b0011100110;
    pxcRom[12477] <= 10'b0100000000;
    pxcRom[12478] <= 10'b0100011111;
    pxcRom[12479] <= 10'b0101001100;
    pxcRom[12480] <= 10'b0101111101;
    pxcRom[12481] <= 10'b0110011001;
    pxcRom[12482] <= 10'b0110010010;
    pxcRom[12483] <= 10'b0110110011;
    pxcRom[12484] <= 10'b0111001101;
    pxcRom[12485] <= 10'b1000100110;
    pxcRom[12486] <= 10'b1000100110;
    pxcRom[12487] <= 10'b1000100110;
    pxcRom[12488] <= 10'b1000100110;
    pxcRom[12489] <= 10'b1000100110;
    pxcRom[12490] <= 10'b1000100110;
    pxcRom[12491] <= 10'b1000100110;
    pxcRom[12492] <= 10'b1000100110;
    pxcRom[12493] <= 10'b1000100110;
    pxcRom[12494] <= 10'b0111111001;
    pxcRom[12495] <= 10'b0111011111;
    pxcRom[12496] <= 10'b0110101001;
    pxcRom[12497] <= 10'b0110000111;
    pxcRom[12498] <= 10'b0101100011;
    pxcRom[12499] <= 10'b0101010011;
    pxcRom[12500] <= 10'b0101010011;
    pxcRom[12501] <= 10'b0101010101;
    pxcRom[12502] <= 10'b0101101001;
    pxcRom[12503] <= 10'b0101100110;
    pxcRom[12504] <= 10'b0101110000;
    pxcRom[12505] <= 10'b0101111000;
    pxcRom[12506] <= 10'b0110010010;
    pxcRom[12507] <= 10'b0110110011;
    pxcRom[12508] <= 10'b0111001101;
    pxcRom[12509] <= 10'b0111011111;
    pxcRom[12510] <= 10'b0111011111;
    pxcRom[12511] <= 10'b1000100110;
    pxcRom[12512] <= 10'b1000100110;
    pxcRom[12513] <= 10'b1000100110;
    pxcRom[12514] <= 10'b1000100110;
    pxcRom[12515] <= 10'b1000100110;
    pxcRom[12516] <= 10'b1000100110;
    pxcRom[12517] <= 10'b1000100110;
    pxcRom[12518] <= 10'b1000100110;
    pxcRom[12519] <= 10'b1000100110;
    pxcRom[12520] <= 10'b1000100110;
    pxcRom[12521] <= 10'b1000100110;
    pxcRom[12522] <= 10'b1000100110;
    pxcRom[12523] <= 10'b1000100110;
    pxcRom[12524] <= 10'b1000100110;
    pxcRom[12525] <= 10'b1000100110;
    pxcRom[12526] <= 10'b0111111001;
    pxcRom[12527] <= 10'b0111111001;
    pxcRom[12528] <= 10'b0111111001;
    pxcRom[12529] <= 10'b0111111001;
    pxcRom[12530] <= 10'b1000100110;
    pxcRom[12531] <= 10'b1000100110;
    pxcRom[12532] <= 10'b1000100110;
    pxcRom[12533] <= 10'b1000100110;
    pxcRom[12534] <= 10'b1000100110;
    pxcRom[12535] <= 10'b1000100110;
    pxcRom[12536] <= 10'b1000100110;
    pxcRom[12537] <= 10'b1000100110;
    pxcRom[12538] <= 10'b1000100110;
    pxcRom[12539] <= 10'b1000100110;
    pxcRom[12540] <= 10'b1000100110;
    pxcRom[12541] <= 10'b1000100110;
    pxcRom[12542] <= 10'b1000100110;
    pxcRom[12543] <= 10'b1000100110;
    pxcRom[12544] <= 10'b1000101011;
    pxcRom[12545] <= 10'b1000101011;
    pxcRom[12546] <= 10'b1000101011;
    pxcRom[12547] <= 10'b1000101011;
    pxcRom[12548] <= 10'b1000101011;
    pxcRom[12549] <= 10'b1000101011;
    pxcRom[12550] <= 10'b1000101011;
    pxcRom[12551] <= 10'b1000101011;
    pxcRom[12552] <= 10'b1000101011;
    pxcRom[12553] <= 10'b1000101011;
    pxcRom[12554] <= 10'b1000101011;
    pxcRom[12555] <= 10'b1000101011;
    pxcRom[12556] <= 10'b0111111111;
    pxcRom[12557] <= 10'b0111111111;
    pxcRom[12558] <= 10'b1000101011;
    pxcRom[12559] <= 10'b1000101011;
    pxcRom[12560] <= 10'b1000101011;
    pxcRom[12561] <= 10'b1000101011;
    pxcRom[12562] <= 10'b1000101011;
    pxcRom[12563] <= 10'b1000101011;
    pxcRom[12564] <= 10'b1000101011;
    pxcRom[12565] <= 10'b1000101011;
    pxcRom[12566] <= 10'b1000101011;
    pxcRom[12567] <= 10'b1000101011;
    pxcRom[12568] <= 10'b1000101011;
    pxcRom[12569] <= 10'b1000101011;
    pxcRom[12570] <= 10'b1000101011;
    pxcRom[12571] <= 10'b1000101011;
    pxcRom[12572] <= 10'b1000101011;
    pxcRom[12573] <= 10'b1000101011;
    pxcRom[12574] <= 10'b1000101011;
    pxcRom[12575] <= 10'b1000101011;
    pxcRom[12576] <= 10'b1000101011;
    pxcRom[12577] <= 10'b0111111111;
    pxcRom[12578] <= 10'b0110111001;
    pxcRom[12579] <= 10'b0110010010;
    pxcRom[12580] <= 10'b0101111110;
    pxcRom[12581] <= 10'b0101100000;
    pxcRom[12582] <= 10'b0101000011;
    pxcRom[12583] <= 10'b0100101001;
    pxcRom[12584] <= 10'b0100100001;
    pxcRom[12585] <= 10'b0100100100;
    pxcRom[12586] <= 10'b0100100010;
    pxcRom[12587] <= 10'b0100101101;
    pxcRom[12588] <= 10'b0100101111;
    pxcRom[12589] <= 10'b0100110100;
    pxcRom[12590] <= 10'b0101000110;
    pxcRom[12591] <= 10'b0101011011;
    pxcRom[12592] <= 10'b0101101100;
    pxcRom[12593] <= 10'b0110011000;
    pxcRom[12594] <= 10'b0111000100;
    pxcRom[12595] <= 10'b0111111111;
    pxcRom[12596] <= 10'b1000101011;
    pxcRom[12597] <= 10'b1000101011;
    pxcRom[12598] <= 10'b1000101011;
    pxcRom[12599] <= 10'b1000101011;
    pxcRom[12600] <= 10'b1000101011;
    pxcRom[12601] <= 10'b1000101011;
    pxcRom[12602] <= 10'b0111111111;
    pxcRom[12603] <= 10'b1000101011;
    pxcRom[12604] <= 10'b0111010011;
    pxcRom[12605] <= 10'b0111010011;
    pxcRom[12606] <= 10'b0101101111;
    pxcRom[12607] <= 10'b0100111000;
    pxcRom[12608] <= 10'b0100011001;
    pxcRom[12609] <= 10'b0011101010;
    pxcRom[12610] <= 10'b0011001011;
    pxcRom[12611] <= 10'b0010101110;
    pxcRom[12612] <= 10'b0010010111;
    pxcRom[12613] <= 10'b0010000010;
    pxcRom[12614] <= 10'b0001110100;
    pxcRom[12615] <= 10'b0001101001;
    pxcRom[12616] <= 10'b0001100111;
    pxcRom[12617] <= 10'b0001101100;
    pxcRom[12618] <= 10'b0001110110;
    pxcRom[12619] <= 10'b0010001010;
    pxcRom[12620] <= 10'b0010101001;
    pxcRom[12621] <= 10'b0011010010;
    pxcRom[12622] <= 10'b0100000000;
    pxcRom[12623] <= 10'b0100111110;
    pxcRom[12624] <= 10'b0110000111;
    pxcRom[12625] <= 10'b0111010011;
    pxcRom[12626] <= 10'b1000101011;
    pxcRom[12627] <= 10'b1000101011;
    pxcRom[12628] <= 10'b1000101011;
    pxcRom[12629] <= 10'b1000101011;
    pxcRom[12630] <= 10'b0111111111;
    pxcRom[12631] <= 10'b0111010011;
    pxcRom[12632] <= 10'b0110111001;
    pxcRom[12633] <= 10'b0110000011;
    pxcRom[12634] <= 10'b0101001100;
    pxcRom[12635] <= 10'b0100010001;
    pxcRom[12636] <= 10'b0011100101;
    pxcRom[12637] <= 10'b0011000000;
    pxcRom[12638] <= 10'b0010011110;
    pxcRom[12639] <= 10'b0010000011;
    pxcRom[12640] <= 10'b0001101011;
    pxcRom[12641] <= 10'b0001010110;
    pxcRom[12642] <= 10'b0001000011;
    pxcRom[12643] <= 10'b0000111000;
    pxcRom[12644] <= 10'b0000110100;
    pxcRom[12645] <= 10'b0000110110;
    pxcRom[12646] <= 10'b0001000000;
    pxcRom[12647] <= 10'b0001010011;
    pxcRom[12648] <= 10'b0001110001;
    pxcRom[12649] <= 10'b0010011010;
    pxcRom[12650] <= 10'b0011000100;
    pxcRom[12651] <= 10'b0100000101;
    pxcRom[12652] <= 10'b0101000011;
    pxcRom[12653] <= 10'b0110011000;
    pxcRom[12654] <= 10'b0111111111;
    pxcRom[12655] <= 10'b1000101011;
    pxcRom[12656] <= 10'b1000101011;
    pxcRom[12657] <= 10'b1000101011;
    pxcRom[12658] <= 10'b1000101011;
    pxcRom[12659] <= 10'b0111010011;
    pxcRom[12660] <= 10'b0110111001;
    pxcRom[12661] <= 10'b0101100000;
    pxcRom[12662] <= 10'b0100100110;
    pxcRom[12663] <= 10'b0011111001;
    pxcRom[12664] <= 10'b0011001001;
    pxcRom[12665] <= 10'b0010100101;
    pxcRom[12666] <= 10'b0010000111;
    pxcRom[12667] <= 10'b0001101101;
    pxcRom[12668] <= 10'b0001010100;
    pxcRom[12669] <= 10'b0001000000;
    pxcRom[12670] <= 10'b0000110001;
    pxcRom[12671] <= 10'b0000101000;
    pxcRom[12672] <= 10'b0000100110;
    pxcRom[12673] <= 10'b0000101100;
    pxcRom[12674] <= 10'b0000111010;
    pxcRom[12675] <= 10'b0001001110;
    pxcRom[12676] <= 10'b0001101110;
    pxcRom[12677] <= 10'b0010010001;
    pxcRom[12678] <= 10'b0010111111;
    pxcRom[12679] <= 10'b0011110111;
    pxcRom[12680] <= 10'b0100110000;
    pxcRom[12681] <= 10'b0101110110;
    pxcRom[12682] <= 10'b0111111111;
    pxcRom[12683] <= 10'b0111111111;
    pxcRom[12684] <= 10'b1000101011;
    pxcRom[12685] <= 10'b1000101011;
    pxcRom[12686] <= 10'b0111000100;
    pxcRom[12687] <= 10'b0111111111;
    pxcRom[12688] <= 10'b0110010010;
    pxcRom[12689] <= 10'b0101010010;
    pxcRom[12690] <= 10'b0100011111;
    pxcRom[12691] <= 10'b0011100010;
    pxcRom[12692] <= 10'b0010110110;
    pxcRom[12693] <= 10'b0010010000;
    pxcRom[12694] <= 10'b0001110100;
    pxcRom[12695] <= 10'b0001011000;
    pxcRom[12696] <= 10'b0001000001;
    pxcRom[12697] <= 10'b0000110000;
    pxcRom[12698] <= 10'b0000100110;
    pxcRom[12699] <= 10'b0000100001;
    pxcRom[12700] <= 10'b0000100101;
    pxcRom[12701] <= 10'b0000110000;
    pxcRom[12702] <= 10'b0001000100;
    pxcRom[12703] <= 10'b0001011110;
    pxcRom[12704] <= 10'b0010000000;
    pxcRom[12705] <= 10'b0010100111;
    pxcRom[12706] <= 10'b0011010010;
    pxcRom[12707] <= 10'b0100000000;
    pxcRom[12708] <= 10'b0100101011;
    pxcRom[12709] <= 10'b0101111010;
    pxcRom[12710] <= 10'b0111100101;
    pxcRom[12711] <= 10'b0111111111;
    pxcRom[12712] <= 10'b1000101011;
    pxcRom[12713] <= 10'b1000101011;
    pxcRom[12714] <= 10'b0111100101;
    pxcRom[12715] <= 10'b1000101011;
    pxcRom[12716] <= 10'b0110011111;
    pxcRom[12717] <= 10'b0101000011;
    pxcRom[12718] <= 10'b0100001001;
    pxcRom[12719] <= 10'b0011001101;
    pxcRom[12720] <= 10'b0010100011;
    pxcRom[12721] <= 10'b0001111110;
    pxcRom[12722] <= 10'b0001100010;
    pxcRom[12723] <= 10'b0001000110;
    pxcRom[12724] <= 10'b0000110011;
    pxcRom[12725] <= 10'b0000100110;
    pxcRom[12726] <= 10'b0000100000;
    pxcRom[12727] <= 10'b0000100010;
    pxcRom[12728] <= 10'b0000101110;
    pxcRom[12729] <= 10'b0001000010;
    pxcRom[12730] <= 10'b0001011100;
    pxcRom[12731] <= 10'b0001111110;
    pxcRom[12732] <= 10'b0010100100;
    pxcRom[12733] <= 10'b0011001010;
    pxcRom[12734] <= 10'b0011110000;
    pxcRom[12735] <= 10'b0100100000;
    pxcRom[12736] <= 10'b0101001100;
    pxcRom[12737] <= 10'b0101111110;
    pxcRom[12738] <= 10'b0111100101;
    pxcRom[12739] <= 10'b0111111111;
    pxcRom[12740] <= 10'b1000101011;
    pxcRom[12741] <= 10'b1000101011;
    pxcRom[12742] <= 10'b1000101011;
    pxcRom[12743] <= 10'b1000101011;
    pxcRom[12744] <= 10'b0110111001;
    pxcRom[12745] <= 10'b0101001100;
    pxcRom[12746] <= 10'b0011111000;
    pxcRom[12747] <= 10'b0010111101;
    pxcRom[12748] <= 10'b0010010000;
    pxcRom[12749] <= 10'b0001101111;
    pxcRom[12750] <= 10'b0001001111;
    pxcRom[12751] <= 10'b0000111000;
    pxcRom[12752] <= 10'b0000101000;
    pxcRom[12753] <= 10'b0000011111;
    pxcRom[12754] <= 10'b0000100000;
    pxcRom[12755] <= 10'b0000101010;
    pxcRom[12756] <= 10'b0000111111;
    pxcRom[12757] <= 10'b0001011011;
    pxcRom[12758] <= 10'b0010000001;
    pxcRom[12759] <= 10'b0010101001;
    pxcRom[12760] <= 10'b0011010000;
    pxcRom[12761] <= 10'b0011101011;
    pxcRom[12762] <= 10'b0100010000;
    pxcRom[12763] <= 10'b0100111001;
    pxcRom[12764] <= 10'b0101100000;
    pxcRom[12765] <= 10'b0110010010;
    pxcRom[12766] <= 10'b0111010011;
    pxcRom[12767] <= 10'b0111111111;
    pxcRom[12768] <= 10'b1000101011;
    pxcRom[12769] <= 10'b1000101011;
    pxcRom[12770] <= 10'b1000101011;
    pxcRom[12771] <= 10'b1000101011;
    pxcRom[12772] <= 10'b0110101111;
    pxcRom[12773] <= 10'b0100111110;
    pxcRom[12774] <= 10'b0011100110;
    pxcRom[12775] <= 10'b0010101001;
    pxcRom[12776] <= 10'b0001111110;
    pxcRom[12777] <= 10'b0001011101;
    pxcRom[12778] <= 10'b0000111111;
    pxcRom[12779] <= 10'b0000101011;
    pxcRom[12780] <= 10'b0000011111;
    pxcRom[12781] <= 10'b0000011100;
    pxcRom[12782] <= 10'b0000100101;
    pxcRom[12783] <= 10'b0000111000;
    pxcRom[12784] <= 10'b0001010111;
    pxcRom[12785] <= 10'b0010000000;
    pxcRom[12786] <= 10'b0010101011;
    pxcRom[12787] <= 10'b0011001111;
    pxcRom[12788] <= 10'b0011011110;
    pxcRom[12789] <= 10'b0011110110;
    pxcRom[12790] <= 10'b0100010001;
    pxcRom[12791] <= 10'b0100111110;
    pxcRom[12792] <= 10'b0101110110;
    pxcRom[12793] <= 10'b0110100110;
    pxcRom[12794] <= 10'b0111010011;
    pxcRom[12795] <= 10'b1000101011;
    pxcRom[12796] <= 10'b1000101011;
    pxcRom[12797] <= 10'b1000101011;
    pxcRom[12798] <= 10'b1000101011;
    pxcRom[12799] <= 10'b1000101011;
    pxcRom[12800] <= 10'b0110100110;
    pxcRom[12801] <= 10'b0100100011;
    pxcRom[12802] <= 10'b0011001110;
    pxcRom[12803] <= 10'b0010010110;
    pxcRom[12804] <= 10'b0001101101;
    pxcRom[12805] <= 10'b0001001100;
    pxcRom[12806] <= 10'b0000110010;
    pxcRom[12807] <= 10'b0000100001;
    pxcRom[12808] <= 10'b0000011010;
    pxcRom[12809] <= 10'b0000011110;
    pxcRom[12810] <= 10'b0000101111;
    pxcRom[12811] <= 10'b0001001110;
    pxcRom[12812] <= 10'b0001110100;
    pxcRom[12813] <= 10'b0010011101;
    pxcRom[12814] <= 10'b0010110011;
    pxcRom[12815] <= 10'b0010111001;
    pxcRom[12816] <= 10'b0010111110;
    pxcRom[12817] <= 10'b0011001101;
    pxcRom[12818] <= 10'b0011101100;
    pxcRom[12819] <= 10'b0100010110;
    pxcRom[12820] <= 10'b0101010100;
    pxcRom[12821] <= 10'b0110011000;
    pxcRom[12822] <= 10'b0111100101;
    pxcRom[12823] <= 10'b1000101011;
    pxcRom[12824] <= 10'b1000101011;
    pxcRom[12825] <= 10'b1000101011;
    pxcRom[12826] <= 10'b1000101011;
    pxcRom[12827] <= 10'b1000101011;
    pxcRom[12828] <= 10'b0110101111;
    pxcRom[12829] <= 10'b0100010001;
    pxcRom[12830] <= 10'b0010111010;
    pxcRom[12831] <= 10'b0010000110;
    pxcRom[12832] <= 10'b0001011101;
    pxcRom[12833] <= 10'b0000111101;
    pxcRom[12834] <= 10'b0000100110;
    pxcRom[12835] <= 10'b0000011001;
    pxcRom[12836] <= 10'b0000011001;
    pxcRom[12837] <= 10'b0000100101;
    pxcRom[12838] <= 10'b0000111111;
    pxcRom[12839] <= 10'b0001100011;
    pxcRom[12840] <= 10'b0010000001;
    pxcRom[12841] <= 10'b0010001010;
    pxcRom[12842] <= 10'b0010000100;
    pxcRom[12843] <= 10'b0010000011;
    pxcRom[12844] <= 10'b0010001000;
    pxcRom[12845] <= 10'b0010011001;
    pxcRom[12846] <= 10'b0010110010;
    pxcRom[12847] <= 10'b0011011111;
    pxcRom[12848] <= 10'b0100011010;
    pxcRom[12849] <= 10'b0110000011;
    pxcRom[12850] <= 10'b0111100101;
    pxcRom[12851] <= 10'b1000101011;
    pxcRom[12852] <= 10'b1000101011;
    pxcRom[12853] <= 10'b1000101011;
    pxcRom[12854] <= 10'b1000101011;
    pxcRom[12855] <= 10'b0111111111;
    pxcRom[12856] <= 10'b0110101111;
    pxcRom[12857] <= 10'b0011111010;
    pxcRom[12858] <= 10'b0010101011;
    pxcRom[12859] <= 10'b0001110111;
    pxcRom[12860] <= 10'b0001001110;
    pxcRom[12861] <= 10'b0000101111;
    pxcRom[12862] <= 10'b0000011100;
    pxcRom[12863] <= 10'b0000010110;
    pxcRom[12864] <= 10'b0000011011;
    pxcRom[12865] <= 10'b0000101110;
    pxcRom[12866] <= 10'b0001001100;
    pxcRom[12867] <= 10'b0001100100;
    pxcRom[12868] <= 10'b0001100010;
    pxcRom[12869] <= 10'b0001011000;
    pxcRom[12870] <= 10'b0001010001;
    pxcRom[12871] <= 10'b0001010011;
    pxcRom[12872] <= 10'b0001011100;
    pxcRom[12873] <= 10'b0001101110;
    pxcRom[12874] <= 10'b0010001001;
    pxcRom[12875] <= 10'b0010101101;
    pxcRom[12876] <= 10'b0011101100;
    pxcRom[12877] <= 10'b0101100000;
    pxcRom[12878] <= 10'b0111010011;
    pxcRom[12879] <= 10'b0111111111;
    pxcRom[12880] <= 10'b1000101011;
    pxcRom[12881] <= 10'b1000101011;
    pxcRom[12882] <= 10'b1000101011;
    pxcRom[12883] <= 10'b0111111111;
    pxcRom[12884] <= 10'b0110101111;
    pxcRom[12885] <= 10'b0011101111;
    pxcRom[12886] <= 10'b0010011101;
    pxcRom[12887] <= 10'b0001101000;
    pxcRom[12888] <= 10'b0001000000;
    pxcRom[12889] <= 10'b0000100100;
    pxcRom[12890] <= 10'b0000010101;
    pxcRom[12891] <= 10'b0000010100;
    pxcRom[12892] <= 10'b0000100001;
    pxcRom[12893] <= 10'b0000110111;
    pxcRom[12894] <= 10'b0001001001;
    pxcRom[12895] <= 10'b0001000101;
    pxcRom[12896] <= 10'b0000111000;
    pxcRom[12897] <= 10'b0000110000;
    pxcRom[12898] <= 10'b0000101110;
    pxcRom[12899] <= 10'b0000110010;
    pxcRom[12900] <= 10'b0000111101;
    pxcRom[12901] <= 10'b0001001110;
    pxcRom[12902] <= 10'b0001100111;
    pxcRom[12903] <= 10'b0010001110;
    pxcRom[12904] <= 10'b0011000010;
    pxcRom[12905] <= 10'b0100110000;
    pxcRom[12906] <= 10'b0111100101;
    pxcRom[12907] <= 10'b0111111111;
    pxcRom[12908] <= 10'b1000101011;
    pxcRom[12909] <= 10'b1000101011;
    pxcRom[12910] <= 10'b1000101011;
    pxcRom[12911] <= 10'b1000101011;
    pxcRom[12912] <= 10'b0110011111;
    pxcRom[12913] <= 10'b0011100101;
    pxcRom[12914] <= 10'b0010001110;
    pxcRom[12915] <= 10'b0001011011;
    pxcRom[12916] <= 10'b0000110011;
    pxcRom[12917] <= 10'b0000011100;
    pxcRom[12918] <= 10'b0000010010;
    pxcRom[12919] <= 10'b0000010110;
    pxcRom[12920] <= 10'b0000100110;
    pxcRom[12921] <= 10'b0000110100;
    pxcRom[12922] <= 10'b0000110010;
    pxcRom[12923] <= 10'b0000100101;
    pxcRom[12924] <= 10'b0000011100;
    pxcRom[12925] <= 10'b0000011001;
    pxcRom[12926] <= 10'b0000011011;
    pxcRom[12927] <= 10'b0000100000;
    pxcRom[12928] <= 10'b0000101010;
    pxcRom[12929] <= 10'b0000111011;
    pxcRom[12930] <= 10'b0001010011;
    pxcRom[12931] <= 10'b0001110110;
    pxcRom[12932] <= 10'b0010100111;
    pxcRom[12933] <= 10'b0100010000;
    pxcRom[12934] <= 10'b0111010011;
    pxcRom[12935] <= 10'b0111111111;
    pxcRom[12936] <= 10'b1000101011;
    pxcRom[12937] <= 10'b1000101011;
    pxcRom[12938] <= 10'b1000101011;
    pxcRom[12939] <= 10'b1000101011;
    pxcRom[12940] <= 10'b0110100110;
    pxcRom[12941] <= 10'b0011010101;
    pxcRom[12942] <= 10'b0010000010;
    pxcRom[12943] <= 10'b0001001101;
    pxcRom[12944] <= 10'b0000101010;
    pxcRom[12945] <= 10'b0000010101;
    pxcRom[12946] <= 10'b0000010000;
    pxcRom[12947] <= 10'b0000011000;
    pxcRom[12948] <= 10'b0000100110;
    pxcRom[12949] <= 10'b0000101000;
    pxcRom[12950] <= 10'b0000011101;
    pxcRom[12951] <= 10'b0000010011;
    pxcRom[12952] <= 10'b0000010001;
    pxcRom[12953] <= 10'b0000010010;
    pxcRom[12954] <= 10'b0000010111;
    pxcRom[12955] <= 10'b0000011011;
    pxcRom[12956] <= 10'b0000100001;
    pxcRom[12957] <= 10'b0000101111;
    pxcRom[12958] <= 10'b0001000111;
    pxcRom[12959] <= 10'b0001101010;
    pxcRom[12960] <= 10'b0010011011;
    pxcRom[12961] <= 10'b0011110110;
    pxcRom[12962] <= 10'b0111010011;
    pxcRom[12963] <= 10'b1000101011;
    pxcRom[12964] <= 10'b1000101011;
    pxcRom[12965] <= 10'b1000101011;
    pxcRom[12966] <= 10'b1000101011;
    pxcRom[12967] <= 10'b1000101011;
    pxcRom[12968] <= 10'b0110010010;
    pxcRom[12969] <= 10'b0011001100;
    pxcRom[12970] <= 10'b0001111000;
    pxcRom[12971] <= 10'b0001000101;
    pxcRom[12972] <= 10'b0000100100;
    pxcRom[12973] <= 10'b0000010010;
    pxcRom[12974] <= 10'b0000001111;
    pxcRom[12975] <= 10'b0000011000;
    pxcRom[12976] <= 10'b0000100001;
    pxcRom[12977] <= 10'b0000011100;
    pxcRom[12978] <= 10'b0000010011;
    pxcRom[12979] <= 10'b0000010001;
    pxcRom[12980] <= 10'b0000010101;
    pxcRom[12981] <= 10'b0000011011;
    pxcRom[12982] <= 10'b0000011100;
    pxcRom[12983] <= 10'b0000011011;
    pxcRom[12984] <= 10'b0000011101;
    pxcRom[12985] <= 10'b0000101010;
    pxcRom[12986] <= 10'b0001000001;
    pxcRom[12987] <= 10'b0001100110;
    pxcRom[12988] <= 10'b0010011001;
    pxcRom[12989] <= 10'b0011101010;
    pxcRom[12990] <= 10'b0110101111;
    pxcRom[12991] <= 10'b1000101011;
    pxcRom[12992] <= 10'b1000101011;
    pxcRom[12993] <= 10'b1000101011;
    pxcRom[12994] <= 10'b1000101011;
    pxcRom[12995] <= 10'b1000101011;
    pxcRom[12996] <= 10'b0101110010;
    pxcRom[12997] <= 10'b0011000011;
    pxcRom[12998] <= 10'b0001110101;
    pxcRom[12999] <= 10'b0001000001;
    pxcRom[13000] <= 10'b0000100000;
    pxcRom[13001] <= 10'b0000010000;
    pxcRom[13002] <= 10'b0000001110;
    pxcRom[13003] <= 10'b0000010110;
    pxcRom[13004] <= 10'b0000011011;
    pxcRom[13005] <= 10'b0000011001;
    pxcRom[13006] <= 10'b0000010110;
    pxcRom[13007] <= 10'b0000011011;
    pxcRom[13008] <= 10'b0000100101;
    pxcRom[13009] <= 10'b0000100111;
    pxcRom[13010] <= 10'b0000011111;
    pxcRom[13011] <= 10'b0000011000;
    pxcRom[13012] <= 10'b0000011011;
    pxcRom[13013] <= 10'b0000101001;
    pxcRom[13014] <= 10'b0001000011;
    pxcRom[13015] <= 10'b0001101101;
    pxcRom[13016] <= 10'b0010011111;
    pxcRom[13017] <= 10'b0011101110;
    pxcRom[13018] <= 10'b0110111001;
    pxcRom[13019] <= 10'b1000101011;
    pxcRom[13020] <= 10'b1000101011;
    pxcRom[13021] <= 10'b1000101011;
    pxcRom[13022] <= 10'b1000101011;
    pxcRom[13023] <= 10'b0111111111;
    pxcRom[13024] <= 10'b0101101001;
    pxcRom[13025] <= 10'b0011000100;
    pxcRom[13026] <= 10'b0001110101;
    pxcRom[13027] <= 10'b0001000001;
    pxcRom[13028] <= 10'b0000100000;
    pxcRom[13029] <= 10'b0000001111;
    pxcRom[13030] <= 10'b0000001100;
    pxcRom[13031] <= 10'b0000010001;
    pxcRom[13032] <= 10'b0000010111;
    pxcRom[13033] <= 10'b0000011001;
    pxcRom[13034] <= 10'b0000011111;
    pxcRom[13035] <= 10'b0000101000;
    pxcRom[13036] <= 10'b0000101100;
    pxcRom[13037] <= 10'b0000100100;
    pxcRom[13038] <= 10'b0000011001;
    pxcRom[13039] <= 10'b0000010011;
    pxcRom[13040] <= 10'b0000011010;
    pxcRom[13041] <= 10'b0000101101;
    pxcRom[13042] <= 10'b0001001100;
    pxcRom[13043] <= 10'b0001111011;
    pxcRom[13044] <= 10'b0010110001;
    pxcRom[13045] <= 10'b0100000011;
    pxcRom[13046] <= 10'b0111010011;
    pxcRom[13047] <= 10'b1000101011;
    pxcRom[13048] <= 10'b1000101011;
    pxcRom[13049] <= 10'b1000101011;
    pxcRom[13050] <= 10'b1000101011;
    pxcRom[13051] <= 10'b0111100101;
    pxcRom[13052] <= 10'b0101011000;
    pxcRom[13053] <= 10'b0011001111;
    pxcRom[13054] <= 10'b0001111110;
    pxcRom[13055] <= 10'b0001000111;
    pxcRom[13056] <= 10'b0000100100;
    pxcRom[13057] <= 10'b0000010000;
    pxcRom[13058] <= 10'b0000001001;
    pxcRom[13059] <= 10'b0000001011;
    pxcRom[13060] <= 10'b0000010010;
    pxcRom[13061] <= 10'b0000011001;
    pxcRom[13062] <= 10'b0000011111;
    pxcRom[13063] <= 10'b0000100000;
    pxcRom[13064] <= 10'b0000011100;
    pxcRom[13065] <= 10'b0000010011;
    pxcRom[13066] <= 10'b0000001110;
    pxcRom[13067] <= 10'b0000010010;
    pxcRom[13068] <= 10'b0000100000;
    pxcRom[13069] <= 10'b0000111011;
    pxcRom[13070] <= 10'b0001100000;
    pxcRom[13071] <= 10'b0010010010;
    pxcRom[13072] <= 10'b0011010110;
    pxcRom[13073] <= 10'b0100101100;
    pxcRom[13074] <= 10'b0111010011;
    pxcRom[13075] <= 10'b1000101011;
    pxcRom[13076] <= 10'b1000101011;
    pxcRom[13077] <= 10'b1000101011;
    pxcRom[13078] <= 10'b1000101011;
    pxcRom[13079] <= 10'b0111111111;
    pxcRom[13080] <= 10'b0101011101;
    pxcRom[13081] <= 10'b0011100111;
    pxcRom[13082] <= 10'b0010010010;
    pxcRom[13083] <= 10'b0001010110;
    pxcRom[13084] <= 10'b0000101110;
    pxcRom[13085] <= 10'b0000010100;
    pxcRom[13086] <= 10'b0000001000;
    pxcRom[13087] <= 10'b0000000110;
    pxcRom[13088] <= 10'b0000001001;
    pxcRom[13089] <= 10'b0000001110;
    pxcRom[13090] <= 10'b0000010000;
    pxcRom[13091] <= 10'b0000001110;
    pxcRom[13092] <= 10'b0000001011;
    pxcRom[13093] <= 10'b0000001001;
    pxcRom[13094] <= 10'b0000001101;
    pxcRom[13095] <= 10'b0000011010;
    pxcRom[13096] <= 10'b0000110001;
    pxcRom[13097] <= 10'b0001010100;
    pxcRom[13098] <= 10'b0010000000;
    pxcRom[13099] <= 10'b0010111001;
    pxcRom[13100] <= 10'b0100000011;
    pxcRom[13101] <= 10'b0101101100;
    pxcRom[13102] <= 10'b0111111111;
    pxcRom[13103] <= 10'b1000101011;
    pxcRom[13104] <= 10'b1000101011;
    pxcRom[13105] <= 10'b1000101011;
    pxcRom[13106] <= 10'b1000101011;
    pxcRom[13107] <= 10'b1000101011;
    pxcRom[13108] <= 10'b0101110010;
    pxcRom[13109] <= 10'b0100001001;
    pxcRom[13110] <= 10'b0010110101;
    pxcRom[13111] <= 10'b0001110011;
    pxcRom[13112] <= 10'b0001000011;
    pxcRom[13113] <= 10'b0000100011;
    pxcRom[13114] <= 10'b0000001110;
    pxcRom[13115] <= 10'b0000000110;
    pxcRom[13116] <= 10'b0000000011;
    pxcRom[13117] <= 10'b0000000100;
    pxcRom[13118] <= 10'b0000000101;
    pxcRom[13119] <= 10'b0000000101;
    pxcRom[13120] <= 10'b0000000111;
    pxcRom[13121] <= 10'b0000001101;
    pxcRom[13122] <= 10'b0000011011;
    pxcRom[13123] <= 10'b0000110010;
    pxcRom[13124] <= 10'b0001010101;
    pxcRom[13125] <= 10'b0010000000;
    pxcRom[13126] <= 10'b0010110110;
    pxcRom[13127] <= 10'b0011111011;
    pxcRom[13128] <= 10'b0101011000;
    pxcRom[13129] <= 10'b0110101111;
    pxcRom[13130] <= 10'b0111111111;
    pxcRom[13131] <= 10'b1000101011;
    pxcRom[13132] <= 10'b1000101011;
    pxcRom[13133] <= 10'b1000101011;
    pxcRom[13134] <= 10'b1000101011;
    pxcRom[13135] <= 10'b1000101011;
    pxcRom[13136] <= 10'b0111000100;
    pxcRom[13137] <= 10'b0101001000;
    pxcRom[13138] <= 10'b0011101011;
    pxcRom[13139] <= 10'b0010100011;
    pxcRom[13140] <= 10'b0001101100;
    pxcRom[13141] <= 10'b0001000001;
    pxcRom[13142] <= 10'b0000100100;
    pxcRom[13143] <= 10'b0000010011;
    pxcRom[13144] <= 10'b0000001010;
    pxcRom[13145] <= 10'b0000001000;
    pxcRom[13146] <= 10'b0000001001;
    pxcRom[13147] <= 10'b0000001101;
    pxcRom[13148] <= 10'b0000010110;
    pxcRom[13149] <= 10'b0000100111;
    pxcRom[13150] <= 10'b0001000000;
    pxcRom[13151] <= 10'b0001100011;
    pxcRom[13152] <= 10'b0010010000;
    pxcRom[13153] <= 10'b0011000110;
    pxcRom[13154] <= 10'b0100000111;
    pxcRom[13155] <= 10'b0101010000;
    pxcRom[13156] <= 10'b0110101111;
    pxcRom[13157] <= 10'b0111000100;
    pxcRom[13158] <= 10'b0111111111;
    pxcRom[13159] <= 10'b1000101011;
    pxcRom[13160] <= 10'b1000101011;
    pxcRom[13161] <= 10'b1000101011;
    pxcRom[13162] <= 10'b1000101011;
    pxcRom[13163] <= 10'b1000101011;
    pxcRom[13164] <= 10'b1000101011;
    pxcRom[13165] <= 10'b0111010011;
    pxcRom[13166] <= 10'b0101100110;
    pxcRom[13167] <= 10'b0100000000;
    pxcRom[13168] <= 10'b0011000011;
    pxcRom[13169] <= 10'b0010010011;
    pxcRom[13170] <= 10'b0001101100;
    pxcRom[13171] <= 10'b0001010010;
    pxcRom[13172] <= 10'b0001000011;
    pxcRom[13173] <= 10'b0000111101;
    pxcRom[13174] <= 10'b0000111111;
    pxcRom[13175] <= 10'b0001001000;
    pxcRom[13176] <= 10'b0001010111;
    pxcRom[13177] <= 10'b0001110001;
    pxcRom[13178] <= 10'b0010010011;
    pxcRom[13179] <= 10'b0010111111;
    pxcRom[13180] <= 10'b0011110100;
    pxcRom[13181] <= 10'b0100101010;
    pxcRom[13182] <= 10'b0101110010;
    pxcRom[13183] <= 10'b0111000100;
    pxcRom[13184] <= 10'b1000101011;
    pxcRom[13185] <= 10'b0111111111;
    pxcRom[13186] <= 10'b0111111111;
    pxcRom[13187] <= 10'b1000101011;
    pxcRom[13188] <= 10'b1000101011;
    pxcRom[13189] <= 10'b1000101011;
    pxcRom[13190] <= 10'b1000101011;
    pxcRom[13191] <= 10'b1000101011;
    pxcRom[13192] <= 10'b1000101011;
    pxcRom[13193] <= 10'b1000101011;
    pxcRom[13194] <= 10'b1000101011;
    pxcRom[13195] <= 10'b0110111001;
    pxcRom[13196] <= 10'b0101100110;
    pxcRom[13197] <= 10'b0100111000;
    pxcRom[13198] <= 10'b0100010010;
    pxcRom[13199] <= 10'b0011101111;
    pxcRom[13200] <= 10'b0011011010;
    pxcRom[13201] <= 10'b0011001111;
    pxcRom[13202] <= 10'b0011010000;
    pxcRom[13203] <= 10'b0011010110;
    pxcRom[13204] <= 10'b0011100101;
    pxcRom[13205] <= 10'b0100000101;
    pxcRom[13206] <= 10'b0100100100;
    pxcRom[13207] <= 10'b0101000100;
    pxcRom[13208] <= 10'b0101101111;
    pxcRom[13209] <= 10'b0110100110;
    pxcRom[13210] <= 10'b0111010011;
    pxcRom[13211] <= 10'b1000101011;
    pxcRom[13212] <= 10'b1000101011;
    pxcRom[13213] <= 10'b1000101011;
    pxcRom[13214] <= 10'b1000101011;
    pxcRom[13215] <= 10'b1000101011;
    pxcRom[13216] <= 10'b1000101011;
    pxcRom[13217] <= 10'b1000101011;
    pxcRom[13218] <= 10'b1000101011;
    pxcRom[13219] <= 10'b1000101011;
    pxcRom[13220] <= 10'b1000101011;
    pxcRom[13221] <= 10'b1000101011;
    pxcRom[13222] <= 10'b1000101011;
    pxcRom[13223] <= 10'b1000101011;
    pxcRom[13224] <= 10'b1000101011;
    pxcRom[13225] <= 10'b1000101011;
    pxcRom[13226] <= 10'b1000101011;
    pxcRom[13227] <= 10'b0111010011;
    pxcRom[13228] <= 10'b0110100110;
    pxcRom[13229] <= 10'b0110100110;
    pxcRom[13230] <= 10'b0110011111;
    pxcRom[13231] <= 10'b0110001100;
    pxcRom[13232] <= 10'b0110010010;
    pxcRom[13233] <= 10'b0110101111;
    pxcRom[13234] <= 10'b0111000100;
    pxcRom[13235] <= 10'b0111111111;
    pxcRom[13236] <= 10'b0111111111;
    pxcRom[13237] <= 10'b1000101011;
    pxcRom[13238] <= 10'b1000101011;
    pxcRom[13239] <= 10'b1000101011;
    pxcRom[13240] <= 10'b1000101011;
    pxcRom[13241] <= 10'b1000101011;
    pxcRom[13242] <= 10'b1000101011;
    pxcRom[13243] <= 10'b1000101011;
    pxcRom[13244] <= 10'b1000101011;
    pxcRom[13245] <= 10'b1000101011;
    pxcRom[13246] <= 10'b1000101011;
    pxcRom[13247] <= 10'b1000101011;
    pxcRom[13248] <= 10'b1000101011;
    pxcRom[13249] <= 10'b1000101011;
    pxcRom[13250] <= 10'b1000101011;
    pxcRom[13251] <= 10'b1000101011;
    pxcRom[13252] <= 10'b1000101011;
    pxcRom[13253] <= 10'b1000101011;
    pxcRom[13254] <= 10'b1000101011;
    pxcRom[13255] <= 10'b0111111111;
    pxcRom[13256] <= 10'b0111111111;
    pxcRom[13257] <= 10'b1000101011;
    pxcRom[13258] <= 10'b1000101011;
    pxcRom[13259] <= 10'b1000101011;
    pxcRom[13260] <= 10'b1000101011;
    pxcRom[13261] <= 10'b1000101011;
    pxcRom[13262] <= 10'b1000101011;
    pxcRom[13263] <= 10'b1000101011;
    pxcRom[13264] <= 10'b1000101011;
    pxcRom[13265] <= 10'b1000101011;
    pxcRom[13266] <= 10'b1000101011;
    pxcRom[13267] <= 10'b1000101011;
    pxcRom[13268] <= 10'b1000101011;
    pxcRom[13269] <= 10'b1000101011;
    pxcRom[13270] <= 10'b1000101011;
    pxcRom[13271] <= 10'b1000101011;
    pxcRom[13272] <= 10'b1000101011;
    pxcRom[13273] <= 10'b1000101011;
    pxcRom[13274] <= 10'b1000101011;
    pxcRom[13275] <= 10'b1000101011;
    pxcRom[13276] <= 10'b1000101011;
    pxcRom[13277] <= 10'b1000101011;
    pxcRom[13278] <= 10'b1000101011;
    pxcRom[13279] <= 10'b1000101011;
    pxcRom[13280] <= 10'b1000101011;
    pxcRom[13281] <= 10'b1000101011;
    pxcRom[13282] <= 10'b1000101011;
    pxcRom[13283] <= 10'b1000101011;
    pxcRom[13284] <= 10'b1000101011;
    pxcRom[13285] <= 10'b1000101011;
    pxcRom[13286] <= 10'b1000101011;
    pxcRom[13287] <= 10'b1000101011;
    pxcRom[13288] <= 10'b1000101011;
    pxcRom[13289] <= 10'b1000101011;
    pxcRom[13290] <= 10'b1000101011;
    pxcRom[13291] <= 10'b1000101011;
    pxcRom[13292] <= 10'b1000101011;
    pxcRom[13293] <= 10'b1000101011;
    pxcRom[13294] <= 10'b1000101011;
    pxcRom[13295] <= 10'b1000101011;
    pxcRom[13296] <= 10'b1000101011;
    pxcRom[13297] <= 10'b1000101011;
    pxcRom[13298] <= 10'b1000101011;
    pxcRom[13299] <= 10'b1000101011;
    pxcRom[13300] <= 10'b1000101011;
    pxcRom[13301] <= 10'b1000101011;
    pxcRom[13302] <= 10'b1000101011;
    pxcRom[13303] <= 10'b1000101011;
    pxcRom[13304] <= 10'b1000101011;
    pxcRom[13305] <= 10'b1000101011;
    pxcRom[13306] <= 10'b1000101011;
    pxcRom[13307] <= 10'b1000101011;
    pxcRom[13308] <= 10'b1000101011;
    pxcRom[13309] <= 10'b1000101011;
    pxcRom[13310] <= 10'b1000101011;
    pxcRom[13311] <= 10'b1000101011;
    pxcRom[13312] <= 10'b1000101011;
    pxcRom[13313] <= 10'b1000101011;
    pxcRom[13314] <= 10'b1000101011;
    pxcRom[13315] <= 10'b1000101011;
    pxcRom[13316] <= 10'b1000101011;
    pxcRom[13317] <= 10'b1000101011;
    pxcRom[13318] <= 10'b1000101011;
    pxcRom[13319] <= 10'b1000101011;
    pxcRom[13320] <= 10'b1000101011;
    pxcRom[13321] <= 10'b1000101011;
    pxcRom[13322] <= 10'b1000101011;
    pxcRom[13323] <= 10'b1000101011;
    pxcRom[13324] <= 10'b1000101011;
    pxcRom[13325] <= 10'b1000101011;
    pxcRom[13326] <= 10'b1000101011;
    pxcRom[13327] <= 10'b1000101011;
    pxcRom[13328] <= 10'b1000101111;
    pxcRom[13329] <= 10'b1000101111;
    pxcRom[13330] <= 10'b1000101111;
    pxcRom[13331] <= 10'b1000101111;
    pxcRom[13332] <= 10'b1000101111;
    pxcRom[13333] <= 10'b1000101111;
    pxcRom[13334] <= 10'b1000101111;
    pxcRom[13335] <= 10'b1000101111;
    pxcRom[13336] <= 10'b1000101111;
    pxcRom[13337] <= 10'b1000101111;
    pxcRom[13338] <= 10'b1000101111;
    pxcRom[13339] <= 10'b1000101111;
    pxcRom[13340] <= 10'b1000101111;
    pxcRom[13341] <= 10'b1000101111;
    pxcRom[13342] <= 10'b1000101111;
    pxcRom[13343] <= 10'b1000101111;
    pxcRom[13344] <= 10'b1000101111;
    pxcRom[13345] <= 10'b1000101111;
    pxcRom[13346] <= 10'b1000101111;
    pxcRom[13347] <= 10'b1000101111;
    pxcRom[13348] <= 10'b1000101111;
    pxcRom[13349] <= 10'b1000101111;
    pxcRom[13350] <= 10'b1000101111;
    pxcRom[13351] <= 10'b1000101111;
    pxcRom[13352] <= 10'b1000101111;
    pxcRom[13353] <= 10'b1000101111;
    pxcRom[13354] <= 10'b1000101111;
    pxcRom[13355] <= 10'b1000101111;
    pxcRom[13356] <= 10'b1000101111;
    pxcRom[13357] <= 10'b1000101111;
    pxcRom[13358] <= 10'b1000101111;
    pxcRom[13359] <= 10'b1000101111;
    pxcRom[13360] <= 10'b1000101111;
    pxcRom[13361] <= 10'b1000101111;
    pxcRom[13362] <= 10'b1000101111;
    pxcRom[13363] <= 10'b1000101111;
    pxcRom[13364] <= 10'b1000101111;
    pxcRom[13365] <= 10'b1000101111;
    pxcRom[13366] <= 10'b1000101111;
    pxcRom[13367] <= 10'b1000101111;
    pxcRom[13368] <= 10'b1000101111;
    pxcRom[13369] <= 10'b1000101111;
    pxcRom[13370] <= 10'b1000101111;
    pxcRom[13371] <= 10'b1000101111;
    pxcRom[13372] <= 10'b1000101111;
    pxcRom[13373] <= 10'b1000101111;
    pxcRom[13374] <= 10'b1000101111;
    pxcRom[13375] <= 10'b1000101111;
    pxcRom[13376] <= 10'b1000101111;
    pxcRom[13377] <= 10'b1000101111;
    pxcRom[13378] <= 10'b1000101111;
    pxcRom[13379] <= 10'b1000101111;
    pxcRom[13380] <= 10'b1000101111;
    pxcRom[13381] <= 10'b1000101111;
    pxcRom[13382] <= 10'b1000101111;
    pxcRom[13383] <= 10'b1000101111;
    pxcRom[13384] <= 10'b1000101111;
    pxcRom[13385] <= 10'b1000101111;
    pxcRom[13386] <= 10'b1000101111;
    pxcRom[13387] <= 10'b1000101111;
    pxcRom[13388] <= 10'b1000101111;
    pxcRom[13389] <= 10'b1000101111;
    pxcRom[13390] <= 10'b1000101111;
    pxcRom[13391] <= 10'b1000101111;
    pxcRom[13392] <= 10'b1000101111;
    pxcRom[13393] <= 10'b1000101111;
    pxcRom[13394] <= 10'b1000101111;
    pxcRom[13395] <= 10'b1000101111;
    pxcRom[13396] <= 10'b1000101111;
    pxcRom[13397] <= 10'b1000101111;
    pxcRom[13398] <= 10'b1000101111;
    pxcRom[13399] <= 10'b1000101111;
    pxcRom[13400] <= 10'b1000101111;
    pxcRom[13401] <= 10'b1000101111;
    pxcRom[13402] <= 10'b1000101111;
    pxcRom[13403] <= 10'b1000101111;
    pxcRom[13404] <= 10'b1000101111;
    pxcRom[13405] <= 10'b1000101111;
    pxcRom[13406] <= 10'b1000101111;
    pxcRom[13407] <= 10'b1000101111;
    pxcRom[13408] <= 10'b1000101111;
    pxcRom[13409] <= 10'b1000101111;
    pxcRom[13410] <= 10'b1000101111;
    pxcRom[13411] <= 10'b1000101111;
    pxcRom[13412] <= 10'b1000101111;
    pxcRom[13413] <= 10'b1000101111;
    pxcRom[13414] <= 10'b1000101111;
    pxcRom[13415] <= 10'b1000101111;
    pxcRom[13416] <= 10'b1000101111;
    pxcRom[13417] <= 10'b1000101111;
    pxcRom[13418] <= 10'b1000101111;
    pxcRom[13419] <= 10'b1000101111;
    pxcRom[13420] <= 10'b1000101111;
    pxcRom[13421] <= 10'b1000101111;
    pxcRom[13422] <= 10'b1000101111;
    pxcRom[13423] <= 10'b1000101111;
    pxcRom[13424] <= 10'b1000101111;
    pxcRom[13425] <= 10'b1000101111;
    pxcRom[13426] <= 10'b1000101111;
    pxcRom[13427] <= 10'b1000101111;
    pxcRom[13428] <= 10'b1000101111;
    pxcRom[13429] <= 10'b1000101111;
    pxcRom[13430] <= 10'b1000101111;
    pxcRom[13431] <= 10'b1000101111;
    pxcRom[13432] <= 10'b1000101111;
    pxcRom[13433] <= 10'b1000101111;
    pxcRom[13434] <= 10'b1000101111;
    pxcRom[13435] <= 10'b1000101111;
    pxcRom[13436] <= 10'b1000101111;
    pxcRom[13437] <= 10'b1000101111;
    pxcRom[13438] <= 10'b1000101111;
    pxcRom[13439] <= 10'b1000101111;
    pxcRom[13440] <= 10'b1000101111;
    pxcRom[13441] <= 10'b1000101111;
    pxcRom[13442] <= 10'b1000101111;
    pxcRom[13443] <= 10'b1000000011;
    pxcRom[13444] <= 10'b1000000011;
    pxcRom[13445] <= 10'b1000000011;
    pxcRom[13446] <= 10'b1000101111;
    pxcRom[13447] <= 10'b1000000011;
    pxcRom[13448] <= 10'b1000000011;
    pxcRom[13449] <= 10'b1000000011;
    pxcRom[13450] <= 10'b1000101111;
    pxcRom[13451] <= 10'b0111010110;
    pxcRom[13452] <= 10'b0111010110;
    pxcRom[13453] <= 10'b0111010110;
    pxcRom[13454] <= 10'b0111010110;
    pxcRom[13455] <= 10'b0111101001;
    pxcRom[13456] <= 10'b0111101001;
    pxcRom[13457] <= 10'b1000101111;
    pxcRom[13458] <= 10'b1000101111;
    pxcRom[13459] <= 10'b1000101111;
    pxcRom[13460] <= 10'b1000101111;
    pxcRom[13461] <= 10'b1000000011;
    pxcRom[13462] <= 10'b1000000011;
    pxcRom[13463] <= 10'b1000101111;
    pxcRom[13464] <= 10'b1000101111;
    pxcRom[13465] <= 10'b1000101111;
    pxcRom[13466] <= 10'b1000101111;
    pxcRom[13467] <= 10'b1000101111;
    pxcRom[13468] <= 10'b1000101111;
    pxcRom[13469] <= 10'b1000101111;
    pxcRom[13470] <= 10'b1000101111;
    pxcRom[13471] <= 10'b1000000011;
    pxcRom[13472] <= 10'b0111010110;
    pxcRom[13473] <= 10'b0110001011;
    pxcRom[13474] <= 10'b0101100100;
    pxcRom[13475] <= 10'b0100111101;
    pxcRom[13476] <= 10'b0100100110;
    pxcRom[13477] <= 10'b0100011000;
    pxcRom[13478] <= 10'b0100010001;
    pxcRom[13479] <= 10'b0100010001;
    pxcRom[13480] <= 10'b0100001010;
    pxcRom[13481] <= 10'b0100001110;
    pxcRom[13482] <= 10'b0100010010;
    pxcRom[13483] <= 10'b0100010111;
    pxcRom[13484] <= 10'b0100100001;
    pxcRom[13485] <= 10'b0100110101;
    pxcRom[13486] <= 10'b0101010001;
    pxcRom[13487] <= 10'b0101101111;
    pxcRom[13488] <= 10'b0110100010;
    pxcRom[13489] <= 10'b0110111100;
    pxcRom[13490] <= 10'b0111001000;
    pxcRom[13491] <= 10'b1000101111;
    pxcRom[13492] <= 10'b1000101111;
    pxcRom[13493] <= 10'b1000101111;
    pxcRom[13494] <= 10'b1000101111;
    pxcRom[13495] <= 10'b1000101111;
    pxcRom[13496] <= 10'b1000101111;
    pxcRom[13497] <= 10'b1000101111;
    pxcRom[13498] <= 10'b0110100010;
    pxcRom[13499] <= 10'b0110000110;
    pxcRom[13500] <= 10'b0100110011;
    pxcRom[13501] <= 10'b0011110010;
    pxcRom[13502] <= 10'b0011010010;
    pxcRom[13503] <= 10'b0010110101;
    pxcRom[13504] <= 10'b0010011111;
    pxcRom[13505] <= 10'b0010001101;
    pxcRom[13506] <= 10'b0010000001;
    pxcRom[13507] <= 10'b0001111001;
    pxcRom[13508] <= 10'b0001110101;
    pxcRom[13509] <= 10'b0001110011;
    pxcRom[13510] <= 10'b0001110001;
    pxcRom[13511] <= 10'b0001110011;
    pxcRom[13512] <= 10'b0001110101;
    pxcRom[13513] <= 10'b0001111011;
    pxcRom[13514] <= 10'b0010001000;
    pxcRom[13515] <= 10'b0010011000;
    pxcRom[13516] <= 10'b0010110101;
    pxcRom[13517] <= 10'b0011010101;
    pxcRom[13518] <= 10'b0011111110;
    pxcRom[13519] <= 10'b0100111101;
    pxcRom[13520] <= 10'b0110101010;
    pxcRom[13521] <= 10'b1000101111;
    pxcRom[13522] <= 10'b1000101111;
    pxcRom[13523] <= 10'b1000101111;
    pxcRom[13524] <= 10'b1000000011;
    pxcRom[13525] <= 10'b0110101010;
    pxcRom[13526] <= 10'b0101000011;
    pxcRom[13527] <= 10'b0011111101;
    pxcRom[13528] <= 10'b0011000001;
    pxcRom[13529] <= 10'b0010010011;
    pxcRom[13530] <= 10'b0001110101;
    pxcRom[13531] <= 10'b0001011100;
    pxcRom[13532] <= 10'b0001001001;
    pxcRom[13533] <= 10'b0000111011;
    pxcRom[13534] <= 10'b0000110001;
    pxcRom[13535] <= 10'b0000101010;
    pxcRom[13536] <= 10'b0000100110;
    pxcRom[13537] <= 10'b0000100011;
    pxcRom[13538] <= 10'b0000100001;
    pxcRom[13539] <= 10'b0000100001;
    pxcRom[13540] <= 10'b0000100000;
    pxcRom[13541] <= 10'b0000100011;
    pxcRom[13542] <= 10'b0000101001;
    pxcRom[13543] <= 10'b0000110111;
    pxcRom[13544] <= 10'b0001001011;
    pxcRom[13545] <= 10'b0001101011;
    pxcRom[13546] <= 10'b0010010110;
    pxcRom[13547] <= 10'b0011001101;
    pxcRom[13548] <= 10'b0100101100;
    pxcRom[13549] <= 10'b0110010110;
    pxcRom[13550] <= 10'b1000101111;
    pxcRom[13551] <= 10'b1000101111;
    pxcRom[13552] <= 10'b1000000011;
    pxcRom[13553] <= 10'b0101101111;
    pxcRom[13554] <= 10'b0011111100;
    pxcRom[13555] <= 10'b0010111001;
    pxcRom[13556] <= 10'b0010001100;
    pxcRom[13557] <= 10'b0001101001;
    pxcRom[13558] <= 10'b0001001100;
    pxcRom[13559] <= 10'b0000110110;
    pxcRom[13560] <= 10'b0000100111;
    pxcRom[13561] <= 10'b0000011011;
    pxcRom[13562] <= 10'b0000010011;
    pxcRom[13563] <= 10'b0000001110;
    pxcRom[13564] <= 10'b0000001011;
    pxcRom[13565] <= 10'b0000001011;
    pxcRom[13566] <= 10'b0000001010;
    pxcRom[13567] <= 10'b0000001001;
    pxcRom[13568] <= 10'b0000001010;
    pxcRom[13569] <= 10'b0000001011;
    pxcRom[13570] <= 10'b0000010000;
    pxcRom[13571] <= 10'b0000011011;
    pxcRom[13572] <= 10'b0000101111;
    pxcRom[13573] <= 10'b0001001110;
    pxcRom[13574] <= 10'b0001111000;
    pxcRom[13575] <= 10'b0010110000;
    pxcRom[13576] <= 10'b0100000011;
    pxcRom[13577] <= 10'b0110000010;
    pxcRom[13578] <= 10'b1000101111;
    pxcRom[13579] <= 10'b1000101111;
    pxcRom[13580] <= 10'b0111101001;
    pxcRom[13581] <= 10'b0101010101;
    pxcRom[13582] <= 10'b0011100001;
    pxcRom[13583] <= 10'b0010100111;
    pxcRom[13584] <= 10'b0001111100;
    pxcRom[13585] <= 10'b0001011001;
    pxcRom[13586] <= 10'b0001000000;
    pxcRom[13587] <= 10'b0000101100;
    pxcRom[13588] <= 10'b0000011100;
    pxcRom[13589] <= 10'b0000010011;
    pxcRom[13590] <= 10'b0000001101;
    pxcRom[13591] <= 10'b0000001010;
    pxcRom[13592] <= 10'b0000001010;
    pxcRom[13593] <= 10'b0000001011;
    pxcRom[13594] <= 10'b0000001011;
    pxcRom[13595] <= 10'b0000001010;
    pxcRom[13596] <= 10'b0000001000;
    pxcRom[13597] <= 10'b0000000111;
    pxcRom[13598] <= 10'b0000001010;
    pxcRom[13599] <= 10'b0000010011;
    pxcRom[13600] <= 10'b0000100110;
    pxcRom[13601] <= 10'b0001000101;
    pxcRom[13602] <= 10'b0001101111;
    pxcRom[13603] <= 10'b0010101010;
    pxcRom[13604] <= 10'b0100001010;
    pxcRom[13605] <= 10'b0110000010;
    pxcRom[13606] <= 10'b1000000011;
    pxcRom[13607] <= 10'b1000000011;
    pxcRom[13608] <= 10'b0111101001;
    pxcRom[13609] <= 10'b0101001101;
    pxcRom[13610] <= 10'b0011100000;
    pxcRom[13611] <= 10'b0010100110;
    pxcRom[13612] <= 10'b0001111101;
    pxcRom[13613] <= 10'b0001011100;
    pxcRom[13614] <= 10'b0001000010;
    pxcRom[13615] <= 10'b0000101111;
    pxcRom[13616] <= 10'b0000100001;
    pxcRom[13617] <= 10'b0000011001;
    pxcRom[13618] <= 10'b0000010111;
    pxcRom[13619] <= 10'b0000011000;
    pxcRom[13620] <= 10'b0000011100;
    pxcRom[13621] <= 10'b0000100000;
    pxcRom[13622] <= 10'b0000100001;
    pxcRom[13623] <= 10'b0000011101;
    pxcRom[13624] <= 10'b0000010100;
    pxcRom[13625] <= 10'b0000001100;
    pxcRom[13626] <= 10'b0000001010;
    pxcRom[13627] <= 10'b0000010010;
    pxcRom[13628] <= 10'b0000100110;
    pxcRom[13629] <= 10'b0001000111;
    pxcRom[13630] <= 10'b0001110110;
    pxcRom[13631] <= 10'b0010111100;
    pxcRom[13632] <= 10'b0100101010;
    pxcRom[13633] <= 10'b0110001011;
    pxcRom[13634] <= 10'b1000000011;
    pxcRom[13635] <= 10'b1000000011;
    pxcRom[13636] <= 10'b0111010110;
    pxcRom[13637] <= 10'b0101011000;
    pxcRom[13638] <= 10'b0011110000;
    pxcRom[13639] <= 10'b0010110110;
    pxcRom[13640] <= 10'b0010001100;
    pxcRom[13641] <= 10'b0001101101;
    pxcRom[13642] <= 10'b0001010001;
    pxcRom[13643] <= 10'b0000111101;
    pxcRom[13644] <= 10'b0000110000;
    pxcRom[13645] <= 10'b0000101011;
    pxcRom[13646] <= 10'b0000101101;
    pxcRom[13647] <= 10'b0000110101;
    pxcRom[13648] <= 10'b0001000010;
    pxcRom[13649] <= 10'b0001001100;
    pxcRom[13650] <= 10'b0001001101;
    pxcRom[13651] <= 10'b0000111101;
    pxcRom[13652] <= 10'b0000100011;
    pxcRom[13653] <= 10'b0000010000;
    pxcRom[13654] <= 10'b0000001011;
    pxcRom[13655] <= 10'b0000010101;
    pxcRom[13656] <= 10'b0000101100;
    pxcRom[13657] <= 10'b0001010011;
    pxcRom[13658] <= 10'b0010000111;
    pxcRom[13659] <= 10'b0011010110;
    pxcRom[13660] <= 10'b0101001101;
    pxcRom[13661] <= 10'b0111101001;
    pxcRom[13662] <= 10'b1000101111;
    pxcRom[13663] <= 10'b1000101111;
    pxcRom[13664] <= 10'b0111101001;
    pxcRom[13665] <= 10'b0101101111;
    pxcRom[13666] <= 10'b0100010010;
    pxcRom[13667] <= 10'b0011010110;
    pxcRom[13668] <= 10'b0010100101;
    pxcRom[13669] <= 10'b0010000010;
    pxcRom[13670] <= 10'b0001100101;
    pxcRom[13671] <= 10'b0001010000;
    pxcRom[13672] <= 10'b0001000100;
    pxcRom[13673] <= 10'b0001000011;
    pxcRom[13674] <= 10'b0001001011;
    pxcRom[13675] <= 10'b0001011111;
    pxcRom[13676] <= 10'b0001111001;
    pxcRom[13677] <= 10'b0010001001;
    pxcRom[13678] <= 10'b0001111011;
    pxcRom[13679] <= 10'b0001001101;
    pxcRom[13680] <= 10'b0000100011;
    pxcRom[13681] <= 10'b0000001110;
    pxcRom[13682] <= 10'b0000001100;
    pxcRom[13683] <= 10'b0000011010;
    pxcRom[13684] <= 10'b0000110110;
    pxcRom[13685] <= 10'b0001100111;
    pxcRom[13686] <= 10'b0010100010;
    pxcRom[13687] <= 10'b0011111011;
    pxcRom[13688] <= 10'b0101101111;
    pxcRom[13689] <= 10'b0110111100;
    pxcRom[13690] <= 10'b1000000011;
    pxcRom[13691] <= 10'b1000000011;
    pxcRom[13692] <= 10'b1000101111;
    pxcRom[13693] <= 10'b0110101010;
    pxcRom[13694] <= 10'b0101000001;
    pxcRom[13695] <= 10'b0011111001;
    pxcRom[13696] <= 10'b0011000010;
    pxcRom[13697] <= 10'b0010011001;
    pxcRom[13698] <= 10'b0001111110;
    pxcRom[13699] <= 10'b0001100101;
    pxcRom[13700] <= 10'b0001011010;
    pxcRom[13701] <= 10'b0001011100;
    pxcRom[13702] <= 10'b0001101100;
    pxcRom[13703] <= 10'b0010001011;
    pxcRom[13704] <= 10'b0010110100;
    pxcRom[13705] <= 10'b0010110111;
    pxcRom[13706] <= 10'b0010000000;
    pxcRom[13707] <= 10'b0001000000;
    pxcRom[13708] <= 10'b0000011001;
    pxcRom[13709] <= 10'b0000001011;
    pxcRom[13710] <= 10'b0000001110;
    pxcRom[13711] <= 10'b0000100001;
    pxcRom[13712] <= 10'b0001000101;
    pxcRom[13713] <= 10'b0001111011;
    pxcRom[13714] <= 10'b0010111110;
    pxcRom[13715] <= 10'b0100000111;
    pxcRom[13716] <= 10'b0101010011;
    pxcRom[13717] <= 10'b0110100010;
    pxcRom[13718] <= 10'b1000000011;
    pxcRom[13719] <= 10'b1000101111;
    pxcRom[13720] <= 10'b1000101111;
    pxcRom[13721] <= 10'b1000000011;
    pxcRom[13722] <= 10'b0101100110;
    pxcRom[13723] <= 10'b0100100000;
    pxcRom[13724] <= 10'b0011011001;
    pxcRom[13725] <= 10'b0010110010;
    pxcRom[13726] <= 10'b0010010010;
    pxcRom[13727] <= 10'b0001111011;
    pxcRom[13728] <= 10'b0001110011;
    pxcRom[13729] <= 10'b0001111001;
    pxcRom[13730] <= 10'b0010001011;
    pxcRom[13731] <= 10'b0010101010;
    pxcRom[13732] <= 10'b0010111001;
    pxcRom[13733] <= 10'b0010100100;
    pxcRom[13734] <= 10'b0001100010;
    pxcRom[13735] <= 10'b0000101011;
    pxcRom[13736] <= 10'b0000010000;
    pxcRom[13737] <= 10'b0000001010;
    pxcRom[13738] <= 10'b0000010001;
    pxcRom[13739] <= 10'b0000101100;
    pxcRom[13740] <= 10'b0001010111;
    pxcRom[13741] <= 10'b0010001100;
    pxcRom[13742] <= 10'b0011000011;
    pxcRom[13743] <= 10'b0011111001;
    pxcRom[13744] <= 10'b0100110010;
    pxcRom[13745] <= 10'b0110001011;
    pxcRom[13746] <= 10'b1000101111;
    pxcRom[13747] <= 10'b1000101111;
    pxcRom[13748] <= 10'b1000101111;
    pxcRom[13749] <= 10'b1000101111;
    pxcRom[13750] <= 10'b0110101010;
    pxcRom[13751] <= 10'b0101000101;
    pxcRom[13752] <= 10'b0011111001;
    pxcRom[13753] <= 10'b0011001000;
    pxcRom[13754] <= 10'b0010101000;
    pxcRom[13755] <= 10'b0010010011;
    pxcRom[13756] <= 10'b0010001011;
    pxcRom[13757] <= 10'b0010001110;
    pxcRom[13758] <= 10'b0010011001;
    pxcRom[13759] <= 10'b0010100000;
    pxcRom[13760] <= 10'b0010011011;
    pxcRom[13761] <= 10'b0001110111;
    pxcRom[13762] <= 10'b0001000000;
    pxcRom[13763] <= 10'b0000011010;
    pxcRom[13764] <= 10'b0000001011;
    pxcRom[13765] <= 10'b0000001010;
    pxcRom[13766] <= 10'b0000011001;
    pxcRom[13767] <= 10'b0000111010;
    pxcRom[13768] <= 10'b0001100110;
    pxcRom[13769] <= 10'b0010010111;
    pxcRom[13770] <= 10'b0011000100;
    pxcRom[13771] <= 10'b0011110001;
    pxcRom[13772] <= 10'b0100101100;
    pxcRom[13773] <= 10'b0110010110;
    pxcRom[13774] <= 10'b1000101111;
    pxcRom[13775] <= 10'b1000101111;
    pxcRom[13776] <= 10'b1000000011;
    pxcRom[13777] <= 10'b1000101111;
    pxcRom[13778] <= 10'b0111101001;
    pxcRom[13779] <= 10'b0101101100;
    pxcRom[13780] <= 10'b0100010110;
    pxcRom[13781] <= 10'b0011100011;
    pxcRom[13782] <= 10'b0011000000;
    pxcRom[13783] <= 10'b0010101110;
    pxcRom[13784] <= 10'b0010100000;
    pxcRom[13785] <= 10'b0010011100;
    pxcRom[13786] <= 10'b0010011001;
    pxcRom[13787] <= 10'b0010010010;
    pxcRom[13788] <= 10'b0001111111;
    pxcRom[13789] <= 10'b0001010011;
    pxcRom[13790] <= 10'b0000101000;
    pxcRom[13791] <= 10'b0000010001;
    pxcRom[13792] <= 10'b0000001001;
    pxcRom[13793] <= 10'b0000010000;
    pxcRom[13794] <= 10'b0000100111;
    pxcRom[13795] <= 10'b0001001101;
    pxcRom[13796] <= 10'b0001111011;
    pxcRom[13797] <= 10'b0010101000;
    pxcRom[13798] <= 10'b0011010001;
    pxcRom[13799] <= 10'b0011111101;
    pxcRom[13800] <= 10'b0100111110;
    pxcRom[13801] <= 10'b0110111100;
    pxcRom[13802] <= 10'b1000101111;
    pxcRom[13803] <= 10'b1000101111;
    pxcRom[13804] <= 10'b1000101111;
    pxcRom[13805] <= 10'b1000000011;
    pxcRom[13806] <= 10'b1000101111;
    pxcRom[13807] <= 10'b0110010000;
    pxcRom[13808] <= 10'b0100110111;
    pxcRom[13809] <= 10'b0100000110;
    pxcRom[13810] <= 10'b0011100101;
    pxcRom[13811] <= 10'b0011001011;
    pxcRom[13812] <= 10'b0010111001;
    pxcRom[13813] <= 10'b0010101011;
    pxcRom[13814] <= 10'b0010011111;
    pxcRom[13815] <= 10'b0010001000;
    pxcRom[13816] <= 10'b0001100111;
    pxcRom[13817] <= 10'b0000111001;
    pxcRom[13818] <= 10'b0000011011;
    pxcRom[13819] <= 10'b0000001101;
    pxcRom[13820] <= 10'b0000001100;
    pxcRom[13821] <= 10'b0000011100;
    pxcRom[13822] <= 10'b0000111010;
    pxcRom[13823] <= 10'b0001100100;
    pxcRom[13824] <= 10'b0010010110;
    pxcRom[13825] <= 10'b0011000101;
    pxcRom[13826] <= 10'b0011101000;
    pxcRom[13827] <= 10'b0100011011;
    pxcRom[13828] <= 10'b0101000110;
    pxcRom[13829] <= 10'b0110011100;
    pxcRom[13830] <= 10'b0111101001;
    pxcRom[13831] <= 10'b1000101111;
    pxcRom[13832] <= 10'b1000000011;
    pxcRom[13833] <= 10'b1000000011;
    pxcRom[13834] <= 10'b0110111100;
    pxcRom[13835] <= 10'b0110100010;
    pxcRom[13836] <= 10'b0101011111;
    pxcRom[13837] <= 10'b0100101111;
    pxcRom[13838] <= 10'b0100010100;
    pxcRom[13839] <= 10'b0011110001;
    pxcRom[13840] <= 10'b0011011001;
    pxcRom[13841] <= 10'b0011000010;
    pxcRom[13842] <= 10'b0010100101;
    pxcRom[13843] <= 10'b0001111111;
    pxcRom[13844] <= 10'b0001010000;
    pxcRom[13845] <= 10'b0000101001;
    pxcRom[13846] <= 10'b0000010100;
    pxcRom[13847] <= 10'b0000001101;
    pxcRom[13848] <= 10'b0000010100;
    pxcRom[13849] <= 10'b0000101100;
    pxcRom[13850] <= 10'b0001010000;
    pxcRom[13851] <= 10'b0010000001;
    pxcRom[13852] <= 10'b0010110001;
    pxcRom[13853] <= 10'b0011100101;
    pxcRom[13854] <= 10'b0100010000;
    pxcRom[13855] <= 10'b0101000001;
    pxcRom[13856] <= 10'b0101100110;
    pxcRom[13857] <= 10'b0110111100;
    pxcRom[13858] <= 10'b0111101001;
    pxcRom[13859] <= 10'b1000101111;
    pxcRom[13860] <= 10'b1000101111;
    pxcRom[13861] <= 10'b0111010110;
    pxcRom[13862] <= 10'b0111001000;
    pxcRom[13863] <= 10'b0111001000;
    pxcRom[13864] <= 10'b0110001011;
    pxcRom[13865] <= 10'b0101100001;
    pxcRom[13866] <= 10'b0101000101;
    pxcRom[13867] <= 10'b0100011010;
    pxcRom[13868] <= 10'b0011111000;
    pxcRom[13869] <= 10'b0011001100;
    pxcRom[13870] <= 10'b0010011100;
    pxcRom[13871] <= 10'b0001100111;
    pxcRom[13872] <= 10'b0000111100;
    pxcRom[13873] <= 10'b0000100000;
    pxcRom[13874] <= 10'b0000010010;
    pxcRom[13875] <= 10'b0000010010;
    pxcRom[13876] <= 10'b0000100001;
    pxcRom[13877] <= 10'b0000111111;
    pxcRom[13878] <= 10'b0001101000;
    pxcRom[13879] <= 10'b0010011101;
    pxcRom[13880] <= 10'b0011010011;
    pxcRom[13881] <= 10'b0100001101;
    pxcRom[13882] <= 10'b0101000110;
    pxcRom[13883] <= 10'b0110001011;
    pxcRom[13884] <= 10'b0110011100;
    pxcRom[13885] <= 10'b0111010110;
    pxcRom[13886] <= 10'b1000101111;
    pxcRom[13887] <= 10'b1000101111;
    pxcRom[13888] <= 10'b1000101111;
    pxcRom[13889] <= 10'b1000000011;
    pxcRom[13890] <= 10'b1000101111;
    pxcRom[13891] <= 10'b1000000011;
    pxcRom[13892] <= 10'b0110111100;
    pxcRom[13893] <= 10'b0110000010;
    pxcRom[13894] <= 10'b0101101001;
    pxcRom[13895] <= 10'b0100101011;
    pxcRom[13896] <= 10'b0011110000;
    pxcRom[13897] <= 10'b0010110011;
    pxcRom[13898] <= 10'b0001111100;
    pxcRom[13899] <= 10'b0001001111;
    pxcRom[13900] <= 10'b0000101110;
    pxcRom[13901] <= 10'b0000011011;
    pxcRom[13902] <= 10'b0000010100;
    pxcRom[13903] <= 10'b0000011011;
    pxcRom[13904] <= 10'b0000110001;
    pxcRom[13905] <= 10'b0001010001;
    pxcRom[13906] <= 10'b0001111100;
    pxcRom[13907] <= 10'b0010110011;
    pxcRom[13908] <= 10'b0011110001;
    pxcRom[13909] <= 10'b0100110000;
    pxcRom[13910] <= 10'b0101011111;
    pxcRom[13911] <= 10'b0110101010;
    pxcRom[13912] <= 10'b0110111100;
    pxcRom[13913] <= 10'b0111010110;
    pxcRom[13914] <= 10'b1000101111;
    pxcRom[13915] <= 10'b1000101111;
    pxcRom[13916] <= 10'b1000101111;
    pxcRom[13917] <= 10'b1000101111;
    pxcRom[13918] <= 10'b1000101111;
    pxcRom[13919] <= 10'b1000101111;
    pxcRom[13920] <= 10'b0110111100;
    pxcRom[13921] <= 10'b0101101111;
    pxcRom[13922] <= 10'b0100111010;
    pxcRom[13923] <= 10'b0100000110;
    pxcRom[13924] <= 10'b0011000100;
    pxcRom[13925] <= 10'b0010001100;
    pxcRom[13926] <= 10'b0001100001;
    pxcRom[13927] <= 10'b0000111110;
    pxcRom[13928] <= 10'b0000100110;
    pxcRom[13929] <= 10'b0000011010;
    pxcRom[13930] <= 10'b0000011010;
    pxcRom[13931] <= 10'b0000100111;
    pxcRom[13932] <= 10'b0000111110;
    pxcRom[13933] <= 10'b0001100000;
    pxcRom[13934] <= 10'b0010001100;
    pxcRom[13935] <= 10'b0011000100;
    pxcRom[13936] <= 10'b0011111100;
    pxcRom[13937] <= 10'b0100110000;
    pxcRom[13938] <= 10'b0101101001;
    pxcRom[13939] <= 10'b0110101010;
    pxcRom[13940] <= 10'b0110111100;
    pxcRom[13941] <= 10'b0111101001;
    pxcRom[13942] <= 10'b1000101111;
    pxcRom[13943] <= 10'b1000101111;
    pxcRom[13944] <= 10'b1000101111;
    pxcRom[13945] <= 10'b1000101111;
    pxcRom[13946] <= 10'b1000101111;
    pxcRom[13947] <= 10'b0111101001;
    pxcRom[13948] <= 10'b0110001011;
    pxcRom[13949] <= 10'b0101000000;
    pxcRom[13950] <= 10'b0100001111;
    pxcRom[13951] <= 10'b0011001111;
    pxcRom[13952] <= 10'b0010011010;
    pxcRom[13953] <= 10'b0001101110;
    pxcRom[13954] <= 10'b0001001100;
    pxcRom[13955] <= 10'b0000110011;
    pxcRom[13956] <= 10'b0000100011;
    pxcRom[13957] <= 10'b0000011110;
    pxcRom[13958] <= 10'b0000100010;
    pxcRom[13959] <= 10'b0000110010;
    pxcRom[13960] <= 10'b0001001001;
    pxcRom[13961] <= 10'b0001101011;
    pxcRom[13962] <= 10'b0010011000;
    pxcRom[13963] <= 10'b0011001101;
    pxcRom[13964] <= 10'b0100000001;
    pxcRom[13965] <= 10'b0100111010;
    pxcRom[13966] <= 10'b0101101111;
    pxcRom[13967] <= 10'b0111001000;
    pxcRom[13968] <= 10'b0111001000;
    pxcRom[13969] <= 10'b0111101001;
    pxcRom[13970] <= 10'b1000101111;
    pxcRom[13971] <= 10'b1000101111;
    pxcRom[13972] <= 10'b1000101111;
    pxcRom[13973] <= 10'b1000101111;
    pxcRom[13974] <= 10'b1000101111;
    pxcRom[13975] <= 10'b0111101001;
    pxcRom[13976] <= 10'b0101010101;
    pxcRom[13977] <= 10'b0100011000;
    pxcRom[13978] <= 10'b0011011110;
    pxcRom[13979] <= 10'b0010101001;
    pxcRom[13980] <= 10'b0001111111;
    pxcRom[13981] <= 10'b0001011100;
    pxcRom[13982] <= 10'b0001000000;
    pxcRom[13983] <= 10'b0000101101;
    pxcRom[13984] <= 10'b0000100100;
    pxcRom[13985] <= 10'b0000100100;
    pxcRom[13986] <= 10'b0000101011;
    pxcRom[13987] <= 10'b0000111100;
    pxcRom[13988] <= 10'b0001010011;
    pxcRom[13989] <= 10'b0001110011;
    pxcRom[13990] <= 10'b0010011110;
    pxcRom[13991] <= 10'b0011010000;
    pxcRom[13992] <= 10'b0100000101;
    pxcRom[13993] <= 10'b0101000011;
    pxcRom[13994] <= 10'b0101111010;
    pxcRom[13995] <= 10'b0111010110;
    pxcRom[13996] <= 10'b0111001000;
    pxcRom[13997] <= 10'b1000000011;
    pxcRom[13998] <= 10'b1000101111;
    pxcRom[13999] <= 10'b1000101111;
    pxcRom[14000] <= 10'b1000101111;
    pxcRom[14001] <= 10'b1000101111;
    pxcRom[14002] <= 10'b1000000011;
    pxcRom[14003] <= 10'b0110110011;
    pxcRom[14004] <= 10'b0101000001;
    pxcRom[14005] <= 10'b0011111111;
    pxcRom[14006] <= 10'b0011000101;
    pxcRom[14007] <= 10'b0010010101;
    pxcRom[14008] <= 10'b0001110000;
    pxcRom[14009] <= 10'b0001010010;
    pxcRom[14010] <= 10'b0000111011;
    pxcRom[14011] <= 10'b0000101111;
    pxcRom[14012] <= 10'b0000101010;
    pxcRom[14013] <= 10'b0000101100;
    pxcRom[14014] <= 10'b0000110110;
    pxcRom[14015] <= 10'b0001000101;
    pxcRom[14016] <= 10'b0001011011;
    pxcRom[14017] <= 10'b0001111100;
    pxcRom[14018] <= 10'b0010100100;
    pxcRom[14019] <= 10'b0011010100;
    pxcRom[14020] <= 10'b0100000101;
    pxcRom[14021] <= 10'b0101001000;
    pxcRom[14022] <= 10'b0110010000;
    pxcRom[14023] <= 10'b1000000011;
    pxcRom[14024] <= 10'b0111010110;
    pxcRom[14025] <= 10'b1000000011;
    pxcRom[14026] <= 10'b1000101111;
    pxcRom[14027] <= 10'b1000101111;
    pxcRom[14028] <= 10'b1000101111;
    pxcRom[14029] <= 10'b1000101111;
    pxcRom[14030] <= 10'b1000101111;
    pxcRom[14031] <= 10'b0110110011;
    pxcRom[14032] <= 10'b0101011010;
    pxcRom[14033] <= 10'b0100000011;
    pxcRom[14034] <= 10'b0011000100;
    pxcRom[14035] <= 10'b0010010010;
    pxcRom[14036] <= 10'b0001101101;
    pxcRom[14037] <= 10'b0001010011;
    pxcRom[14038] <= 10'b0001000000;
    pxcRom[14039] <= 10'b0000110111;
    pxcRom[14040] <= 10'b0000110101;
    pxcRom[14041] <= 10'b0000111001;
    pxcRom[14042] <= 10'b0001000010;
    pxcRom[14043] <= 10'b0001010011;
    pxcRom[14044] <= 10'b0001101000;
    pxcRom[14045] <= 10'b0010000111;
    pxcRom[14046] <= 10'b0010110000;
    pxcRom[14047] <= 10'b0011010111;
    pxcRom[14048] <= 10'b0100001100;
    pxcRom[14049] <= 10'b0101001100;
    pxcRom[14050] <= 10'b0101111010;
    pxcRom[14051] <= 10'b0111010110;
    pxcRom[14052] <= 10'b0111010110;
    pxcRom[14053] <= 10'b1000101111;
    pxcRom[14054] <= 10'b1000101111;
    pxcRom[14055] <= 10'b1000101111;
    pxcRom[14056] <= 10'b1000101111;
    pxcRom[14057] <= 10'b1000101111;
    pxcRom[14058] <= 10'b1000101111;
    pxcRom[14059] <= 10'b1000101111;
    pxcRom[14060] <= 10'b0110010000;
    pxcRom[14061] <= 10'b0100110001;
    pxcRom[14062] <= 10'b0011101011;
    pxcRom[14063] <= 10'b0010110011;
    pxcRom[14064] <= 10'b0010010000;
    pxcRom[14065] <= 10'b0001110111;
    pxcRom[14066] <= 10'b0001100101;
    pxcRom[14067] <= 10'b0001011010;
    pxcRom[14068] <= 10'b0001010111;
    pxcRom[14069] <= 10'b0001011001;
    pxcRom[14070] <= 10'b0001100010;
    pxcRom[14071] <= 10'b0001110001;
    pxcRom[14072] <= 10'b0010000101;
    pxcRom[14073] <= 10'b0010100010;
    pxcRom[14074] <= 10'b0011000101;
    pxcRom[14075] <= 10'b0011110001;
    pxcRom[14076] <= 10'b0100110011;
    pxcRom[14077] <= 10'b0101011100;
    pxcRom[14078] <= 10'b0110001011;
    pxcRom[14079] <= 10'b0111010110;
    pxcRom[14080] <= 10'b1000101111;
    pxcRom[14081] <= 10'b1000000011;
    pxcRom[14082] <= 10'b1000101111;
    pxcRom[14083] <= 10'b1000101111;
    pxcRom[14084] <= 10'b1000101111;
    pxcRom[14085] <= 10'b1000101111;
    pxcRom[14086] <= 10'b1000101111;
    pxcRom[14087] <= 10'b1000101111;
    pxcRom[14088] <= 10'b0111101001;
    pxcRom[14089] <= 10'b0110110011;
    pxcRom[14090] <= 10'b0101110011;
    pxcRom[14091] <= 10'b0101001101;
    pxcRom[14092] <= 10'b0100110000;
    pxcRom[14093] <= 10'b0100011110;
    pxcRom[14094] <= 10'b0011111000;
    pxcRom[14095] <= 10'b0011101111;
    pxcRom[14096] <= 10'b0011100000;
    pxcRom[14097] <= 10'b0011010110;
    pxcRom[14098] <= 10'b0011010010;
    pxcRom[14099] <= 10'b0011011010;
    pxcRom[14100] <= 10'b0011100101;
    pxcRom[14101] <= 10'b0011111100;
    pxcRom[14102] <= 10'b0100011100;
    pxcRom[14103] <= 10'b0101001111;
    pxcRom[14104] <= 10'b0110010110;
    pxcRom[14105] <= 10'b0110110011;
    pxcRom[14106] <= 10'b0111001000;
    pxcRom[14107] <= 10'b0111101001;
    pxcRom[14108] <= 10'b1000101111;
    pxcRom[14109] <= 10'b1000101111;
    pxcRom[14110] <= 10'b1000101111;
    pxcRom[14111] <= 10'b1000101111;
    pxcRom[14112] <= 10'b1000101011;
    pxcRom[14113] <= 10'b1000101011;
    pxcRom[14114] <= 10'b1000101011;
    pxcRom[14115] <= 10'b1000101011;
    pxcRom[14116] <= 10'b1000101011;
    pxcRom[14117] <= 10'b1000101011;
    pxcRom[14118] <= 10'b1000101011;
    pxcRom[14119] <= 10'b1000101011;
    pxcRom[14120] <= 10'b1000101011;
    pxcRom[14121] <= 10'b1000101011;
    pxcRom[14122] <= 10'b1000101011;
    pxcRom[14123] <= 10'b1000101011;
    pxcRom[14124] <= 10'b1000101011;
    pxcRom[14125] <= 10'b1000101011;
    pxcRom[14126] <= 10'b1000101011;
    pxcRom[14127] <= 10'b1000101011;
    pxcRom[14128] <= 10'b1000101011;
    pxcRom[14129] <= 10'b1000101011;
    pxcRom[14130] <= 10'b1000101011;
    pxcRom[14131] <= 10'b1000101011;
    pxcRom[14132] <= 10'b1000101011;
    pxcRom[14133] <= 10'b1000101011;
    pxcRom[14134] <= 10'b1000101011;
    pxcRom[14135] <= 10'b1000101011;
    pxcRom[14136] <= 10'b1000101011;
    pxcRom[14137] <= 10'b1000101011;
    pxcRom[14138] <= 10'b1000101011;
    pxcRom[14139] <= 10'b1000101011;
    pxcRom[14140] <= 10'b1000101011;
    pxcRom[14141] <= 10'b1000101011;
    pxcRom[14142] <= 10'b1000101011;
    pxcRom[14143] <= 10'b1000101011;
    pxcRom[14144] <= 10'b1000101011;
    pxcRom[14145] <= 10'b1000101011;
    pxcRom[14146] <= 10'b1000101011;
    pxcRom[14147] <= 10'b1000101011;
    pxcRom[14148] <= 10'b1000101011;
    pxcRom[14149] <= 10'b1000101011;
    pxcRom[14150] <= 10'b1000101011;
    pxcRom[14151] <= 10'b1000101011;
    pxcRom[14152] <= 10'b1000101011;
    pxcRom[14153] <= 10'b1000101011;
    pxcRom[14154] <= 10'b1000101011;
    pxcRom[14155] <= 10'b1000101011;
    pxcRom[14156] <= 10'b1000101011;
    pxcRom[14157] <= 10'b1000101011;
    pxcRom[14158] <= 10'b1000101011;
    pxcRom[14159] <= 10'b1000101011;
    pxcRom[14160] <= 10'b1000101011;
    pxcRom[14161] <= 10'b1000101011;
    pxcRom[14162] <= 10'b1000101011;
    pxcRom[14163] <= 10'b1000101011;
    pxcRom[14164] <= 10'b1000101011;
    pxcRom[14165] <= 10'b1000101011;
    pxcRom[14166] <= 10'b1000101011;
    pxcRom[14167] <= 10'b1000101011;
    pxcRom[14168] <= 10'b1000101011;
    pxcRom[14169] <= 10'b1000101011;
    pxcRom[14170] <= 10'b1000101011;
    pxcRom[14171] <= 10'b1000101011;
    pxcRom[14172] <= 10'b1000101011;
    pxcRom[14173] <= 10'b1000101011;
    pxcRom[14174] <= 10'b1000101011;
    pxcRom[14175] <= 10'b1000101011;
    pxcRom[14176] <= 10'b1000101011;
    pxcRom[14177] <= 10'b1000101011;
    pxcRom[14178] <= 10'b1000101011;
    pxcRom[14179] <= 10'b1000101011;
    pxcRom[14180] <= 10'b1000101011;
    pxcRom[14181] <= 10'b1000101011;
    pxcRom[14182] <= 10'b1000101011;
    pxcRom[14183] <= 10'b1000101011;
    pxcRom[14184] <= 10'b1000101011;
    pxcRom[14185] <= 10'b0111111110;
    pxcRom[14186] <= 10'b0111111110;
    pxcRom[14187] <= 10'b1000101011;
    pxcRom[14188] <= 10'b1000101011;
    pxcRom[14189] <= 10'b1000101011;
    pxcRom[14190] <= 10'b1000101011;
    pxcRom[14191] <= 10'b1000101011;
    pxcRom[14192] <= 10'b1000101011;
    pxcRom[14193] <= 10'b1000101011;
    pxcRom[14194] <= 10'b1000101011;
    pxcRom[14195] <= 10'b1000101011;
    pxcRom[14196] <= 10'b1000101011;
    pxcRom[14197] <= 10'b1000101011;
    pxcRom[14198] <= 10'b1000101011;
    pxcRom[14199] <= 10'b1000101011;
    pxcRom[14200] <= 10'b1000101011;
    pxcRom[14201] <= 10'b1000101011;
    pxcRom[14202] <= 10'b1000101011;
    pxcRom[14203] <= 10'b1000101011;
    pxcRom[14204] <= 10'b0111111110;
    pxcRom[14205] <= 10'b0111111110;
    pxcRom[14206] <= 10'b0111000100;
    pxcRom[14207] <= 10'b0110101110;
    pxcRom[14208] <= 10'b0110010001;
    pxcRom[14209] <= 10'b0101110101;
    pxcRom[14210] <= 10'b0101101011;
    pxcRom[14211] <= 10'b0101011000;
    pxcRom[14212] <= 10'b0101000101;
    pxcRom[14213] <= 10'b0101010101;
    pxcRom[14214] <= 10'b0101010101;
    pxcRom[14215] <= 10'b0101101110;
    pxcRom[14216] <= 10'b0110000111;
    pxcRom[14217] <= 10'b0110010001;
    pxcRom[14218] <= 10'b0110011110;
    pxcRom[14219] <= 10'b0111000100;
    pxcRom[14220] <= 10'b0111100100;
    pxcRom[14221] <= 10'b0111111110;
    pxcRom[14222] <= 10'b1000101011;
    pxcRom[14223] <= 10'b1000101011;
    pxcRom[14224] <= 10'b1000101011;
    pxcRom[14225] <= 10'b1000101011;
    pxcRom[14226] <= 10'b1000101011;
    pxcRom[14227] <= 10'b1000101011;
    pxcRom[14228] <= 10'b1000101011;
    pxcRom[14229] <= 10'b0111111110;
    pxcRom[14230] <= 10'b0111111110;
    pxcRom[14231] <= 10'b0110010111;
    pxcRom[14232] <= 10'b0101000101;
    pxcRom[14233] <= 10'b0100010010;
    pxcRom[14234] <= 10'b0011101000;
    pxcRom[14235] <= 10'b0011000000;
    pxcRom[14236] <= 10'b0010011110;
    pxcRom[14237] <= 10'b0010000100;
    pxcRom[14238] <= 10'b0001110011;
    pxcRom[14239] <= 10'b0001101011;
    pxcRom[14240] <= 10'b0001101011;
    pxcRom[14241] <= 10'b0001110000;
    pxcRom[14242] <= 10'b0001111111;
    pxcRom[14243] <= 10'b0010010110;
    pxcRom[14244] <= 10'b0010101101;
    pxcRom[14245] <= 10'b0011001110;
    pxcRom[14246] <= 10'b0011110110;
    pxcRom[14247] <= 10'b0100110010;
    pxcRom[14248] <= 10'b0101011010;
    pxcRom[14249] <= 10'b0110000111;
    pxcRom[14250] <= 10'b0111000100;
    pxcRom[14251] <= 10'b0111111110;
    pxcRom[14252] <= 10'b1000101011;
    pxcRom[14253] <= 10'b1000101011;
    pxcRom[14254] <= 10'b1000101011;
    pxcRom[14255] <= 10'b1000101011;
    pxcRom[14256] <= 10'b0111111110;
    pxcRom[14257] <= 10'b0110111000;
    pxcRom[14258] <= 10'b0101010101;
    pxcRom[14259] <= 10'b0100010000;
    pxcRom[14260] <= 10'b0011010001;
    pxcRom[14261] <= 10'b0010100001;
    pxcRom[14262] <= 10'b0001111010;
    pxcRom[14263] <= 10'b0001010111;
    pxcRom[14264] <= 10'b0000111100;
    pxcRom[14265] <= 10'b0000101010;
    pxcRom[14266] <= 10'b0000011110;
    pxcRom[14267] <= 10'b0000010111;
    pxcRom[14268] <= 10'b0000010110;
    pxcRom[14269] <= 10'b0000011010;
    pxcRom[14270] <= 10'b0000100101;
    pxcRom[14271] <= 10'b0000110110;
    pxcRom[14272] <= 10'b0001001100;
    pxcRom[14273] <= 10'b0001101001;
    pxcRom[14274] <= 10'b0010001011;
    pxcRom[14275] <= 10'b0010111000;
    pxcRom[14276] <= 10'b0011101000;
    pxcRom[14277] <= 10'b0100100011;
    pxcRom[14278] <= 10'b0101111101;
    pxcRom[14279] <= 10'b0111111110;
    pxcRom[14280] <= 10'b1000101011;
    pxcRom[14281] <= 10'b1000101011;
    pxcRom[14282] <= 10'b1000101011;
    pxcRom[14283] <= 10'b1000101011;
    pxcRom[14284] <= 10'b0110011110;
    pxcRom[14285] <= 10'b0101001111;
    pxcRom[14286] <= 10'b0011111111;
    pxcRom[14287] <= 10'b0010111110;
    pxcRom[14288] <= 10'b0010001111;
    pxcRom[14289] <= 10'b0001100110;
    pxcRom[14290] <= 10'b0001000101;
    pxcRom[14291] <= 10'b0000101100;
    pxcRom[14292] <= 10'b0000011011;
    pxcRom[14293] <= 10'b0000010000;
    pxcRom[14294] <= 10'b0000001011;
    pxcRom[14295] <= 10'b0000001001;
    pxcRom[14296] <= 10'b0000001001;
    pxcRom[14297] <= 10'b0000001100;
    pxcRom[14298] <= 10'b0000010011;
    pxcRom[14299] <= 10'b0000011110;
    pxcRom[14300] <= 10'b0000101111;
    pxcRom[14301] <= 10'b0001000110;
    pxcRom[14302] <= 10'b0001100100;
    pxcRom[14303] <= 10'b0010000111;
    pxcRom[14304] <= 10'b0010110110;
    pxcRom[14305] <= 10'b0011110110;
    pxcRom[14306] <= 10'b0101011010;
    pxcRom[14307] <= 10'b0111100100;
    pxcRom[14308] <= 10'b1000101011;
    pxcRom[14309] <= 10'b1000101011;
    pxcRom[14310] <= 10'b1000101011;
    pxcRom[14311] <= 10'b0111111110;
    pxcRom[14312] <= 10'b0101011010;
    pxcRom[14313] <= 10'b0100001110;
    pxcRom[14314] <= 10'b0011000101;
    pxcRom[14315] <= 10'b0010010000;
    pxcRom[14316] <= 10'b0001101000;
    pxcRom[14317] <= 10'b0001000110;
    pxcRom[14318] <= 10'b0000101100;
    pxcRom[14319] <= 10'b0000011010;
    pxcRom[14320] <= 10'b0000010001;
    pxcRom[14321] <= 10'b0000001101;
    pxcRom[14322] <= 10'b0000001110;
    pxcRom[14323] <= 10'b0000001111;
    pxcRom[14324] <= 10'b0000010001;
    pxcRom[14325] <= 10'b0000010001;
    pxcRom[14326] <= 10'b0000010011;
    pxcRom[14327] <= 10'b0000011000;
    pxcRom[14328] <= 10'b0000100100;
    pxcRom[14329] <= 10'b0000111000;
    pxcRom[14330] <= 10'b0001010000;
    pxcRom[14331] <= 10'b0001101110;
    pxcRom[14332] <= 10'b0010011100;
    pxcRom[14333] <= 10'b0011100010;
    pxcRom[14334] <= 10'b0100110110;
    pxcRom[14335] <= 10'b0111000100;
    pxcRom[14336] <= 10'b1000101011;
    pxcRom[14337] <= 10'b1000101011;
    pxcRom[14338] <= 10'b1000101011;
    pxcRom[14339] <= 10'b0110010111;
    pxcRom[14340] <= 10'b0100110000;
    pxcRom[14341] <= 10'b0011100111;
    pxcRom[14342] <= 10'b0010100110;
    pxcRom[14343] <= 10'b0001111000;
    pxcRom[14344] <= 10'b0001010010;
    pxcRom[14345] <= 10'b0000110100;
    pxcRom[14346] <= 10'b0000100000;
    pxcRom[14347] <= 10'b0000010101;
    pxcRom[14348] <= 10'b0000010011;
    pxcRom[14349] <= 10'b0000010111;
    pxcRom[14350] <= 10'b0000100000;
    pxcRom[14351] <= 10'b0000100111;
    pxcRom[14352] <= 10'b0000100110;
    pxcRom[14353] <= 10'b0000100010;
    pxcRom[14354] <= 10'b0000011011;
    pxcRom[14355] <= 10'b0000011001;
    pxcRom[14356] <= 10'b0000100001;
    pxcRom[14357] <= 10'b0000110001;
    pxcRom[14358] <= 10'b0001000110;
    pxcRom[14359] <= 10'b0001100111;
    pxcRom[14360] <= 10'b0010010000;
    pxcRom[14361] <= 10'b0011010001;
    pxcRom[14362] <= 10'b0100110010;
    pxcRom[14363] <= 10'b0110111000;
    pxcRom[14364] <= 10'b1000101011;
    pxcRom[14365] <= 10'b1000101011;
    pxcRom[14366] <= 10'b1000101011;
    pxcRom[14367] <= 10'b0110010111;
    pxcRom[14368] <= 10'b0100011001;
    pxcRom[14369] <= 10'b0011010110;
    pxcRom[14370] <= 10'b0010010111;
    pxcRom[14371] <= 10'b0001101011;
    pxcRom[14372] <= 10'b0001000111;
    pxcRom[14373] <= 10'b0000101011;
    pxcRom[14374] <= 10'b0000011100;
    pxcRom[14375] <= 10'b0000010111;
    pxcRom[14376] <= 10'b0000011011;
    pxcRom[14377] <= 10'b0000101000;
    pxcRom[14378] <= 10'b0000111010;
    pxcRom[14379] <= 10'b0001000011;
    pxcRom[14380] <= 10'b0000111011;
    pxcRom[14381] <= 10'b0000101010;
    pxcRom[14382] <= 10'b0000011101;
    pxcRom[14383] <= 10'b0000011001;
    pxcRom[14384] <= 10'b0000100000;
    pxcRom[14385] <= 10'b0000110001;
    pxcRom[14386] <= 10'b0001001000;
    pxcRom[14387] <= 10'b0001101001;
    pxcRom[14388] <= 10'b0010010001;
    pxcRom[14389] <= 10'b0011010110;
    pxcRom[14390] <= 10'b0100110011;
    pxcRom[14391] <= 10'b0110111000;
    pxcRom[14392] <= 10'b1000101011;
    pxcRom[14393] <= 10'b1000101011;
    pxcRom[14394] <= 10'b1000101011;
    pxcRom[14395] <= 10'b0110100110;
    pxcRom[14396] <= 10'b0100010101;
    pxcRom[14397] <= 10'b0011001110;
    pxcRom[14398] <= 10'b0010010101;
    pxcRom[14399] <= 10'b0001100111;
    pxcRom[14400] <= 10'b0001000100;
    pxcRom[14401] <= 10'b0000101010;
    pxcRom[14402] <= 10'b0000011100;
    pxcRom[14403] <= 10'b0000011001;
    pxcRom[14404] <= 10'b0000100000;
    pxcRom[14405] <= 10'b0000110011;
    pxcRom[14406] <= 10'b0001000111;
    pxcRom[14407] <= 10'b0001001000;
    pxcRom[14408] <= 10'b0000110110;
    pxcRom[14409] <= 10'b0000100010;
    pxcRom[14410] <= 10'b0000010111;
    pxcRom[14411] <= 10'b0000011000;
    pxcRom[14412] <= 10'b0000100010;
    pxcRom[14413] <= 10'b0000110111;
    pxcRom[14414] <= 10'b0001010011;
    pxcRom[14415] <= 10'b0001111000;
    pxcRom[14416] <= 10'b0010100101;
    pxcRom[14417] <= 10'b0011100011;
    pxcRom[14418] <= 10'b0101001001;
    pxcRom[14419] <= 10'b0110111000;
    pxcRom[14420] <= 10'b1000101011;
    pxcRom[14421] <= 10'b1000101011;
    pxcRom[14422] <= 10'b1000101011;
    pxcRom[14423] <= 10'b0110100110;
    pxcRom[14424] <= 10'b0100011110;
    pxcRom[14425] <= 10'b0011001111;
    pxcRom[14426] <= 10'b0010010111;
    pxcRom[14427] <= 10'b0001101010;
    pxcRom[14428] <= 10'b0001001000;
    pxcRom[14429] <= 10'b0000101101;
    pxcRom[14430] <= 10'b0000011110;
    pxcRom[14431] <= 10'b0000011000;
    pxcRom[14432] <= 10'b0000011101;
    pxcRom[14433] <= 10'b0000101010;
    pxcRom[14434] <= 10'b0000110111;
    pxcRom[14435] <= 10'b0000110001;
    pxcRom[14436] <= 10'b0000100000;
    pxcRom[14437] <= 10'b0000010101;
    pxcRom[14438] <= 10'b0000010011;
    pxcRom[14439] <= 10'b0000011100;
    pxcRom[14440] <= 10'b0000101110;
    pxcRom[14441] <= 10'b0001001001;
    pxcRom[14442] <= 10'b0001101011;
    pxcRom[14443] <= 10'b0010010111;
    pxcRom[14444] <= 10'b0011000101;
    pxcRom[14445] <= 10'b0100000111;
    pxcRom[14446] <= 10'b0101011010;
    pxcRom[14447] <= 10'b0111111110;
    pxcRom[14448] <= 10'b1000101011;
    pxcRom[14449] <= 10'b1000101011;
    pxcRom[14450] <= 10'b1000101011;
    pxcRom[14451] <= 10'b0111000100;
    pxcRom[14452] <= 10'b0100111010;
    pxcRom[14453] <= 10'b0011100010;
    pxcRom[14454] <= 10'b0010100111;
    pxcRom[14455] <= 10'b0001111010;
    pxcRom[14456] <= 10'b0001010010;
    pxcRom[14457] <= 10'b0000110110;
    pxcRom[14458] <= 10'b0000100010;
    pxcRom[14459] <= 10'b0000010111;
    pxcRom[14460] <= 10'b0000010101;
    pxcRom[14461] <= 10'b0000011010;
    pxcRom[14462] <= 10'b0000011111;
    pxcRom[14463] <= 10'b0000010111;
    pxcRom[14464] <= 10'b0000010000;
    pxcRom[14465] <= 10'b0000001111;
    pxcRom[14466] <= 10'b0000010111;
    pxcRom[14467] <= 10'b0000101000;
    pxcRom[14468] <= 10'b0001000100;
    pxcRom[14469] <= 10'b0001100110;
    pxcRom[14470] <= 10'b0010001111;
    pxcRom[14471] <= 10'b0010111101;
    pxcRom[14472] <= 10'b0011101000;
    pxcRom[14473] <= 10'b0100110110;
    pxcRom[14474] <= 10'b0110000010;
    pxcRom[14475] <= 10'b0111100100;
    pxcRom[14476] <= 10'b1000101011;
    pxcRom[14477] <= 10'b1000101011;
    pxcRom[14478] <= 10'b1000101011;
    pxcRom[14479] <= 10'b0111010010;
    pxcRom[14480] <= 10'b0101011010;
    pxcRom[14481] <= 10'b0100000110;
    pxcRom[14482] <= 10'b0011000011;
    pxcRom[14483] <= 10'b0010001111;
    pxcRom[14484] <= 10'b0001100101;
    pxcRom[14485] <= 10'b0001000011;
    pxcRom[14486] <= 10'b0000101010;
    pxcRom[14487] <= 10'b0000010111;
    pxcRom[14488] <= 10'b0000001101;
    pxcRom[14489] <= 10'b0000001100;
    pxcRom[14490] <= 10'b0000001101;
    pxcRom[14491] <= 10'b0000001001;
    pxcRom[14492] <= 10'b0000001001;
    pxcRom[14493] <= 10'b0000010010;
    pxcRom[14494] <= 10'b0000100100;
    pxcRom[14495] <= 10'b0001000001;
    pxcRom[14496] <= 10'b0001100101;
    pxcRom[14497] <= 10'b0010001111;
    pxcRom[14498] <= 10'b0010111001;
    pxcRom[14499] <= 10'b0011101001;
    pxcRom[14500] <= 10'b0100011100;
    pxcRom[14501] <= 10'b0101011111;
    pxcRom[14502] <= 10'b0110111000;
    pxcRom[14503] <= 10'b0111111110;
    pxcRom[14504] <= 10'b1000101011;
    pxcRom[14505] <= 10'b1000101011;
    pxcRom[14506] <= 10'b1000101011;
    pxcRom[14507] <= 10'b0111111110;
    pxcRom[14508] <= 10'b0110010111;
    pxcRom[14509] <= 10'b0100101010;
    pxcRom[14510] <= 10'b0011100110;
    pxcRom[14511] <= 10'b0010101100;
    pxcRom[14512] <= 10'b0001111100;
    pxcRom[14513] <= 10'b0001010100;
    pxcRom[14514] <= 10'b0000110001;
    pxcRom[14515] <= 10'b0000011000;
    pxcRom[14516] <= 10'b0000001010;
    pxcRom[14517] <= 10'b0000000101;
    pxcRom[14518] <= 10'b0000000100;
    pxcRom[14519] <= 10'b0000000101;
    pxcRom[14520] <= 10'b0000001011;
    pxcRom[14521] <= 10'b0000011100;
    pxcRom[14522] <= 10'b0000111010;
    pxcRom[14523] <= 10'b0001011111;
    pxcRom[14524] <= 10'b0010000111;
    pxcRom[14525] <= 10'b0010101101;
    pxcRom[14526] <= 10'b0011010101;
    pxcRom[14527] <= 10'b0100000010;
    pxcRom[14528] <= 10'b0100111010;
    pxcRom[14529] <= 10'b0101110101;
    pxcRom[14530] <= 10'b0111111110;
    pxcRom[14531] <= 10'b1000101011;
    pxcRom[14532] <= 10'b1000101011;
    pxcRom[14533] <= 10'b1000101011;
    pxcRom[14534] <= 10'b1000101011;
    pxcRom[14535] <= 10'b0111111110;
    pxcRom[14536] <= 10'b0111010010;
    pxcRom[14537] <= 10'b0101000111;
    pxcRom[14538] <= 10'b0011111010;
    pxcRom[14539] <= 10'b0010111011;
    pxcRom[14540] <= 10'b0010000110;
    pxcRom[14541] <= 10'b0001011001;
    pxcRom[14542] <= 10'b0000110010;
    pxcRom[14543] <= 10'b0000010110;
    pxcRom[14544] <= 10'b0000001000;
    pxcRom[14545] <= 10'b0000000100;
    pxcRom[14546] <= 10'b0000000101;
    pxcRom[14547] <= 10'b0000001000;
    pxcRom[14548] <= 10'b0000010010;
    pxcRom[14549] <= 10'b0000101010;
    pxcRom[14550] <= 10'b0001001010;
    pxcRom[14551] <= 10'b0001101101;
    pxcRom[14552] <= 10'b0010010000;
    pxcRom[14553] <= 10'b0010110110;
    pxcRom[14554] <= 10'b0011011100;
    pxcRom[14555] <= 10'b0100001001;
    pxcRom[14556] <= 10'b0100111010;
    pxcRom[14557] <= 10'b0110010111;
    pxcRom[14558] <= 10'b1000101011;
    pxcRom[14559] <= 10'b1000101011;
    pxcRom[14560] <= 10'b1000101011;
    pxcRom[14561] <= 10'b1000101011;
    pxcRom[14562] <= 10'b1000101011;
    pxcRom[14563] <= 10'b0111111110;
    pxcRom[14564] <= 10'b0111000100;
    pxcRom[14565] <= 10'b0100111101;
    pxcRom[14566] <= 10'b0011100110;
    pxcRom[14567] <= 10'b0010101001;
    pxcRom[14568] <= 10'b0001110101;
    pxcRom[14569] <= 10'b0001001001;
    pxcRom[14570] <= 10'b0000100111;
    pxcRom[14571] <= 10'b0000010001;
    pxcRom[14572] <= 10'b0000001001;
    pxcRom[14573] <= 10'b0000001001;
    pxcRom[14574] <= 10'b0000001100;
    pxcRom[14575] <= 10'b0000010000;
    pxcRom[14576] <= 10'b0000011100;
    pxcRom[14577] <= 10'b0000101111;
    pxcRom[14578] <= 10'b0001001010;
    pxcRom[14579] <= 10'b0001101001;
    pxcRom[14580] <= 10'b0010001001;
    pxcRom[14581] <= 10'b0010101100;
    pxcRom[14582] <= 10'b0011010010;
    pxcRom[14583] <= 10'b0011111001;
    pxcRom[14584] <= 10'b0100101001;
    pxcRom[14585] <= 10'b0110010111;
    pxcRom[14586] <= 10'b1000101011;
    pxcRom[14587] <= 10'b1000101011;
    pxcRom[14588] <= 10'b1000101011;
    pxcRom[14589] <= 10'b1000101011;
    pxcRom[14590] <= 10'b1000101011;
    pxcRom[14591] <= 10'b0111100100;
    pxcRom[14592] <= 10'b0110000111;
    pxcRom[14593] <= 10'b0100010111;
    pxcRom[14594] <= 10'b0011000100;
    pxcRom[14595] <= 10'b0010001000;
    pxcRom[14596] <= 10'b0001011000;
    pxcRom[14597] <= 10'b0000110011;
    pxcRom[14598] <= 10'b0000011011;
    pxcRom[14599] <= 10'b0000001111;
    pxcRom[14600] <= 10'b0000001110;
    pxcRom[14601] <= 10'b0000010100;
    pxcRom[14602] <= 10'b0000011010;
    pxcRom[14603] <= 10'b0000011100;
    pxcRom[14604] <= 10'b0000100001;
    pxcRom[14605] <= 10'b0000101111;
    pxcRom[14606] <= 10'b0001000100;
    pxcRom[14607] <= 10'b0001011111;
    pxcRom[14608] <= 10'b0001111101;
    pxcRom[14609] <= 10'b0010011111;
    pxcRom[14610] <= 10'b0011000001;
    pxcRom[14611] <= 10'b0011101001;
    pxcRom[14612] <= 10'b0100011111;
    pxcRom[14613] <= 10'b0110101110;
    pxcRom[14614] <= 10'b0111111110;
    pxcRom[14615] <= 10'b1000101011;
    pxcRom[14616] <= 10'b1000101011;
    pxcRom[14617] <= 10'b1000101011;
    pxcRom[14618] <= 10'b1000101011;
    pxcRom[14619] <= 10'b0111111110;
    pxcRom[14620] <= 10'b0101100010;
    pxcRom[14621] <= 10'b0011100111;
    pxcRom[14622] <= 10'b0010100010;
    pxcRom[14623] <= 10'b0001101011;
    pxcRom[14624] <= 10'b0001000000;
    pxcRom[14625] <= 10'b0000100101;
    pxcRom[14626] <= 10'b0000010101;
    pxcRom[14627] <= 10'b0000010010;
    pxcRom[14628] <= 10'b0000011010;
    pxcRom[14629] <= 10'b0000100110;
    pxcRom[14630] <= 10'b0000101010;
    pxcRom[14631] <= 10'b0000100100;
    pxcRom[14632] <= 10'b0000100100;
    pxcRom[14633] <= 10'b0000101110;
    pxcRom[14634] <= 10'b0000111110;
    pxcRom[14635] <= 10'b0001010110;
    pxcRom[14636] <= 10'b0001110010;
    pxcRom[14637] <= 10'b0010010100;
    pxcRom[14638] <= 10'b0010110111;
    pxcRom[14639] <= 10'b0011011110;
    pxcRom[14640] <= 10'b0100100010;
    pxcRom[14641] <= 10'b0110101110;
    pxcRom[14642] <= 10'b0111111110;
    pxcRom[14643] <= 10'b1000101011;
    pxcRom[14644] <= 10'b1000101011;
    pxcRom[14645] <= 10'b1000101011;
    pxcRom[14646] <= 10'b1000101011;
    pxcRom[14647] <= 10'b0111100100;
    pxcRom[14648] <= 10'b0100111000;
    pxcRom[14649] <= 10'b0011000111;
    pxcRom[14650] <= 10'b0010000111;
    pxcRom[14651] <= 10'b0001010101;
    pxcRom[14652] <= 10'b0000110011;
    pxcRom[14653] <= 10'b0000011110;
    pxcRom[14654] <= 10'b0000010110;
    pxcRom[14655] <= 10'b0000011011;
    pxcRom[14656] <= 10'b0000101001;
    pxcRom[14657] <= 10'b0000110110;
    pxcRom[14658] <= 10'b0000110011;
    pxcRom[14659] <= 10'b0000101001;
    pxcRom[14660] <= 10'b0000100101;
    pxcRom[14661] <= 10'b0000101011;
    pxcRom[14662] <= 10'b0000111001;
    pxcRom[14663] <= 10'b0001010001;
    pxcRom[14664] <= 10'b0001101100;
    pxcRom[14665] <= 10'b0010001111;
    pxcRom[14666] <= 10'b0010110101;
    pxcRom[14667] <= 10'b0011100010;
    pxcRom[14668] <= 10'b0100111000;
    pxcRom[14669] <= 10'b0111010010;
    pxcRom[14670] <= 10'b1000101011;
    pxcRom[14671] <= 10'b1000101011;
    pxcRom[14672] <= 10'b1000101011;
    pxcRom[14673] <= 10'b1000101011;
    pxcRom[14674] <= 10'b1000101011;
    pxcRom[14675] <= 10'b0111010010;
    pxcRom[14676] <= 10'b0100100110;
    pxcRom[14677] <= 10'b0010111000;
    pxcRom[14678] <= 10'b0001110101;
    pxcRom[14679] <= 10'b0001001001;
    pxcRom[14680] <= 10'b0000101101;
    pxcRom[14681] <= 10'b0000011101;
    pxcRom[14682] <= 10'b0000011000;
    pxcRom[14683] <= 10'b0000100001;
    pxcRom[14684] <= 10'b0000101101;
    pxcRom[14685] <= 10'b0000110100;
    pxcRom[14686] <= 10'b0000101100;
    pxcRom[14687] <= 10'b0000100101;
    pxcRom[14688] <= 10'b0000100010;
    pxcRom[14689] <= 10'b0000101000;
    pxcRom[14690] <= 10'b0000110111;
    pxcRom[14691] <= 10'b0001001111;
    pxcRom[14692] <= 10'b0001101100;
    pxcRom[14693] <= 10'b0010010001;
    pxcRom[14694] <= 10'b0010111100;
    pxcRom[14695] <= 10'b0011110000;
    pxcRom[14696] <= 10'b0101010101;
    pxcRom[14697] <= 10'b0111010010;
    pxcRom[14698] <= 10'b1000101011;
    pxcRom[14699] <= 10'b1000101011;
    pxcRom[14700] <= 10'b1000101011;
    pxcRom[14701] <= 10'b1000101011;
    pxcRom[14702] <= 10'b1000101011;
    pxcRom[14703] <= 10'b0111010010;
    pxcRom[14704] <= 10'b0100100101;
    pxcRom[14705] <= 10'b0010110011;
    pxcRom[14706] <= 10'b0001110001;
    pxcRom[14707] <= 10'b0001000111;
    pxcRom[14708] <= 10'b0000101101;
    pxcRom[14709] <= 10'b0000011101;
    pxcRom[14710] <= 10'b0000010111;
    pxcRom[14711] <= 10'b0000011000;
    pxcRom[14712] <= 10'b0000011100;
    pxcRom[14713] <= 10'b0000011101;
    pxcRom[14714] <= 10'b0000011011;
    pxcRom[14715] <= 10'b0000011001;
    pxcRom[14716] <= 10'b0000011101;
    pxcRom[14717] <= 10'b0000100111;
    pxcRom[14718] <= 10'b0000111001;
    pxcRom[14719] <= 10'b0001010011;
    pxcRom[14720] <= 10'b0001110101;
    pxcRom[14721] <= 10'b0010011101;
    pxcRom[14722] <= 10'b0011001011;
    pxcRom[14723] <= 10'b0100001000;
    pxcRom[14724] <= 10'b0110000010;
    pxcRom[14725] <= 10'b0111111110;
    pxcRom[14726] <= 10'b1000101011;
    pxcRom[14727] <= 10'b1000101011;
    pxcRom[14728] <= 10'b1000101011;
    pxcRom[14729] <= 10'b1000101011;
    pxcRom[14730] <= 10'b1000101011;
    pxcRom[14731] <= 10'b0111010010;
    pxcRom[14732] <= 10'b0100111010;
    pxcRom[14733] <= 10'b0010111001;
    pxcRom[14734] <= 10'b0001111000;
    pxcRom[14735] <= 10'b0001001111;
    pxcRom[14736] <= 10'b0000110011;
    pxcRom[14737] <= 10'b0000100000;
    pxcRom[14738] <= 10'b0000010011;
    pxcRom[14739] <= 10'b0000001101;
    pxcRom[14740] <= 10'b0000001011;
    pxcRom[14741] <= 10'b0000001011;
    pxcRom[14742] <= 10'b0000001101;
    pxcRom[14743] <= 10'b0000010010;
    pxcRom[14744] <= 10'b0000011100;
    pxcRom[14745] <= 10'b0000101101;
    pxcRom[14746] <= 10'b0001000011;
    pxcRom[14747] <= 10'b0001100011;
    pxcRom[14748] <= 10'b0010001000;
    pxcRom[14749] <= 10'b0010111000;
    pxcRom[14750] <= 10'b0011100111;
    pxcRom[14751] <= 10'b0100110110;
    pxcRom[14752] <= 10'b0110011110;
    pxcRom[14753] <= 10'b0111100100;
    pxcRom[14754] <= 10'b1000101011;
    pxcRom[14755] <= 10'b1000101011;
    pxcRom[14756] <= 10'b1000101011;
    pxcRom[14757] <= 10'b1000101011;
    pxcRom[14758] <= 10'b1000101011;
    pxcRom[14759] <= 10'b0111100100;
    pxcRom[14760] <= 10'b0101101011;
    pxcRom[14761] <= 10'b0011011100;
    pxcRom[14762] <= 10'b0010001110;
    pxcRom[14763] <= 10'b0001100010;
    pxcRom[14764] <= 10'b0001000001;
    pxcRom[14765] <= 10'b0000101011;
    pxcRom[14766] <= 10'b0000011010;
    pxcRom[14767] <= 10'b0000001111;
    pxcRom[14768] <= 10'b0000001010;
    pxcRom[14769] <= 10'b0000001010;
    pxcRom[14770] <= 10'b0000001111;
    pxcRom[14771] <= 10'b0000011001;
    pxcRom[14772] <= 10'b0000101001;
    pxcRom[14773] <= 10'b0000111111;
    pxcRom[14774] <= 10'b0001011101;
    pxcRom[14775] <= 10'b0010000011;
    pxcRom[14776] <= 10'b0010101111;
    pxcRom[14777] <= 10'b0011100001;
    pxcRom[14778] <= 10'b0100010110;
    pxcRom[14779] <= 10'b0101100101;
    pxcRom[14780] <= 10'b0110111000;
    pxcRom[14781] <= 10'b0111111110;
    pxcRom[14782] <= 10'b1000101011;
    pxcRom[14783] <= 10'b1000101011;
    pxcRom[14784] <= 10'b1000101011;
    pxcRom[14785] <= 10'b1000101011;
    pxcRom[14786] <= 10'b1000101011;
    pxcRom[14787] <= 10'b1000101011;
    pxcRom[14788] <= 10'b0111010010;
    pxcRom[14789] <= 10'b0100101110;
    pxcRom[14790] <= 10'b0011001101;
    pxcRom[14791] <= 10'b0010010110;
    pxcRom[14792] <= 10'b0001101100;
    pxcRom[14793] <= 10'b0001010000;
    pxcRom[14794] <= 10'b0000111100;
    pxcRom[14795] <= 10'b0000101111;
    pxcRom[14796] <= 10'b0000101001;
    pxcRom[14797] <= 10'b0000101001;
    pxcRom[14798] <= 10'b0000110010;
    pxcRom[14799] <= 10'b0001000000;
    pxcRom[14800] <= 10'b0001010101;
    pxcRom[14801] <= 10'b0001110010;
    pxcRom[14802] <= 10'b0010011000;
    pxcRom[14803] <= 10'b0011000001;
    pxcRom[14804] <= 10'b0011110001;
    pxcRom[14805] <= 10'b0100101000;
    pxcRom[14806] <= 10'b0101011101;
    pxcRom[14807] <= 10'b0110111000;
    pxcRom[14808] <= 10'b1000101011;
    pxcRom[14809] <= 10'b1000101011;
    pxcRom[14810] <= 10'b1000101011;
    pxcRom[14811] <= 10'b1000101011;
    pxcRom[14812] <= 10'b1000101011;
    pxcRom[14813] <= 10'b1000101011;
    pxcRom[14814] <= 10'b1000101011;
    pxcRom[14815] <= 10'b1000101011;
    pxcRom[14816] <= 10'b1000101011;
    pxcRom[14817] <= 10'b0111000100;
    pxcRom[14818] <= 10'b0101010101;
    pxcRom[14819] <= 10'b0100100111;
    pxcRom[14820] <= 10'b0100000000;
    pxcRom[14821] <= 10'b0011100110;
    pxcRom[14822] <= 10'b0011010000;
    pxcRom[14823] <= 10'b0011000101;
    pxcRom[14824] <= 10'b0010111111;
    pxcRom[14825] <= 10'b0010111010;
    pxcRom[14826] <= 10'b0010111101;
    pxcRom[14827] <= 10'b0011001011;
    pxcRom[14828] <= 10'b0011100001;
    pxcRom[14829] <= 10'b0100000011;
    pxcRom[14830] <= 10'b0100100000;
    pxcRom[14831] <= 10'b0101000000;
    pxcRom[14832] <= 10'b0101111001;
    pxcRom[14833] <= 10'b0111100100;
    pxcRom[14834] <= 10'b0111111110;
    pxcRom[14835] <= 10'b0111111110;
    pxcRom[14836] <= 10'b1000101011;
    pxcRom[14837] <= 10'b1000101011;
    pxcRom[14838] <= 10'b1000101011;
    pxcRom[14839] <= 10'b1000101011;
    pxcRom[14840] <= 10'b1000101011;
    pxcRom[14841] <= 10'b1000101011;
    pxcRom[14842] <= 10'b1000101011;
    pxcRom[14843] <= 10'b1000101011;
    pxcRom[14844] <= 10'b1000101011;
    pxcRom[14845] <= 10'b1000101011;
    pxcRom[14846] <= 10'b1000101011;
    pxcRom[14847] <= 10'b0111111110;
    pxcRom[14848] <= 10'b0111000100;
    pxcRom[14849] <= 10'b0110111000;
    pxcRom[14850] <= 10'b0110111000;
    pxcRom[14851] <= 10'b0110100110;
    pxcRom[14852] <= 10'b0110100110;
    pxcRom[14853] <= 10'b0110111000;
    pxcRom[14854] <= 10'b0111010010;
    pxcRom[14855] <= 10'b0111100100;
    pxcRom[14856] <= 10'b0111111110;
    pxcRom[14857] <= 10'b0111111110;
    pxcRom[14858] <= 10'b0111111110;
    pxcRom[14859] <= 10'b0111111110;
    pxcRom[14860] <= 10'b1000101011;
    pxcRom[14861] <= 10'b1000101011;
    pxcRom[14862] <= 10'b0111111110;
    pxcRom[14863] <= 10'b1000101011;
    pxcRom[14864] <= 10'b1000101011;
    pxcRom[14865] <= 10'b1000101011;
    pxcRom[14866] <= 10'b1000101011;
    pxcRom[14867] <= 10'b1000101011;
    pxcRom[14868] <= 10'b1000101011;
    pxcRom[14869] <= 10'b1000101011;
    pxcRom[14870] <= 10'b1000101011;
    pxcRom[14871] <= 10'b1000101011;
    pxcRom[14872] <= 10'b1000101011;
    pxcRom[14873] <= 10'b1000101011;
    pxcRom[14874] <= 10'b1000101011;
    pxcRom[14875] <= 10'b1000101011;
    pxcRom[14876] <= 10'b1000101011;
    pxcRom[14877] <= 10'b1000101011;
    pxcRom[14878] <= 10'b1000101011;
    pxcRom[14879] <= 10'b1000101011;
    pxcRom[14880] <= 10'b1000101011;
    pxcRom[14881] <= 10'b1000101011;
    pxcRom[14882] <= 10'b1000101011;
    pxcRom[14883] <= 10'b1000101011;
    pxcRom[14884] <= 10'b1000101011;
    pxcRom[14885] <= 10'b1000101011;
    pxcRom[14886] <= 10'b1000101011;
    pxcRom[14887] <= 10'b1000101011;
    pxcRom[14888] <= 10'b1000101011;
    pxcRom[14889] <= 10'b1000101011;
    pxcRom[14890] <= 10'b1000101011;
    pxcRom[14891] <= 10'b1000101011;
    pxcRom[14892] <= 10'b1000101011;
    pxcRom[14893] <= 10'b1000101011;
    pxcRom[14894] <= 10'b1000101011;
    pxcRom[14895] <= 10'b1000101011;
    pxcRom[14896] <= 10'b1000101100;
    pxcRom[14897] <= 10'b1000101100;
    pxcRom[14898] <= 10'b1000101100;
    pxcRom[14899] <= 10'b1000101100;
    pxcRom[14900] <= 10'b1000101100;
    pxcRom[14901] <= 10'b1000101100;
    pxcRom[14902] <= 10'b1000101100;
    pxcRom[14903] <= 10'b1000101100;
    pxcRom[14904] <= 10'b1000101100;
    pxcRom[14905] <= 10'b1000101100;
    pxcRom[14906] <= 10'b1000101100;
    pxcRom[14907] <= 10'b1000101100;
    pxcRom[14908] <= 10'b1000101100;
    pxcRom[14909] <= 10'b1000101100;
    pxcRom[14910] <= 10'b1000101100;
    pxcRom[14911] <= 10'b1000101100;
    pxcRom[14912] <= 10'b1000101100;
    pxcRom[14913] <= 10'b1000101100;
    pxcRom[14914] <= 10'b1000101100;
    pxcRom[14915] <= 10'b1000101100;
    pxcRom[14916] <= 10'b1000101100;
    pxcRom[14917] <= 10'b1000101100;
    pxcRom[14918] <= 10'b1000101100;
    pxcRom[14919] <= 10'b1000101100;
    pxcRom[14920] <= 10'b1000101100;
    pxcRom[14921] <= 10'b1000101100;
    pxcRom[14922] <= 10'b1000101100;
    pxcRom[14923] <= 10'b1000101100;
    pxcRom[14924] <= 10'b1000101100;
    pxcRom[14925] <= 10'b1000101100;
    pxcRom[14926] <= 10'b1000101100;
    pxcRom[14927] <= 10'b1000101100;
    pxcRom[14928] <= 10'b1000101100;
    pxcRom[14929] <= 10'b1000101100;
    pxcRom[14930] <= 10'b1000101100;
    pxcRom[14931] <= 10'b1000101100;
    pxcRom[14932] <= 10'b1000101100;
    pxcRom[14933] <= 10'b1000101100;
    pxcRom[14934] <= 10'b1000101100;
    pxcRom[14935] <= 10'b1000101100;
    pxcRom[14936] <= 10'b1000101100;
    pxcRom[14937] <= 10'b1000101100;
    pxcRom[14938] <= 10'b1000101100;
    pxcRom[14939] <= 10'b1000101100;
    pxcRom[14940] <= 10'b1000101100;
    pxcRom[14941] <= 10'b1000101100;
    pxcRom[14942] <= 10'b1000101100;
    pxcRom[14943] <= 10'b1000101100;
    pxcRom[14944] <= 10'b1000101100;
    pxcRom[14945] <= 10'b1000101100;
    pxcRom[14946] <= 10'b1000101100;
    pxcRom[14947] <= 10'b1000101100;
    pxcRom[14948] <= 10'b1000101100;
    pxcRom[14949] <= 10'b1000101100;
    pxcRom[14950] <= 10'b1000101100;
    pxcRom[14951] <= 10'b1000101100;
    pxcRom[14952] <= 10'b1000101100;
    pxcRom[14953] <= 10'b1000101100;
    pxcRom[14954] <= 10'b1000101100;
    pxcRom[14955] <= 10'b1000101100;
    pxcRom[14956] <= 10'b1000101100;
    pxcRom[14957] <= 10'b1000101100;
    pxcRom[14958] <= 10'b1000101100;
    pxcRom[14959] <= 10'b1000101100;
    pxcRom[14960] <= 10'b1000101100;
    pxcRom[14961] <= 10'b1000101100;
    pxcRom[14962] <= 10'b1000101100;
    pxcRom[14963] <= 10'b1000101100;
    pxcRom[14964] <= 10'b1000101100;
    pxcRom[14965] <= 10'b1000101100;
    pxcRom[14966] <= 10'b1000101100;
    pxcRom[14967] <= 10'b1000101100;
    pxcRom[14968] <= 10'b1000101100;
    pxcRom[14969] <= 10'b1000101100;
    pxcRom[14970] <= 10'b1000101100;
    pxcRom[14971] <= 10'b1000101100;
    pxcRom[14972] <= 10'b1000101100;
    pxcRom[14973] <= 10'b1000101100;
    pxcRom[14974] <= 10'b1000101100;
    pxcRom[14975] <= 10'b1000101100;
    pxcRom[14976] <= 10'b1000101100;
    pxcRom[14977] <= 10'b1000101100;
    pxcRom[14978] <= 10'b1000101100;
    pxcRom[14979] <= 10'b1000101100;
    pxcRom[14980] <= 10'b1000101100;
    pxcRom[14981] <= 10'b1000101100;
    pxcRom[14982] <= 10'b1000101100;
    pxcRom[14983] <= 10'b1000101100;
    pxcRom[14984] <= 10'b1000101100;
    pxcRom[14985] <= 10'b1000101100;
    pxcRom[14986] <= 10'b1000101100;
    pxcRom[14987] <= 10'b1000101100;
    pxcRom[14988] <= 10'b1000101100;
    pxcRom[14989] <= 10'b1000101100;
    pxcRom[14990] <= 10'b1000101100;
    pxcRom[14991] <= 10'b1000101100;
    pxcRom[14992] <= 10'b1000101100;
    pxcRom[14993] <= 10'b1000101100;
    pxcRom[14994] <= 10'b1000101100;
    pxcRom[14995] <= 10'b1000101100;
    pxcRom[14996] <= 10'b1000101100;
    pxcRom[14997] <= 10'b1000101100;
    pxcRom[14998] <= 10'b0111111111;
    pxcRom[14999] <= 10'b1000101100;
    pxcRom[15000] <= 10'b1000101100;
    pxcRom[15001] <= 10'b1000101100;
    pxcRom[15002] <= 10'b1000101100;
    pxcRom[15003] <= 10'b1000101100;
    pxcRom[15004] <= 10'b1000101100;
    pxcRom[15005] <= 10'b1000101100;
    pxcRom[15006] <= 10'b1000101100;
    pxcRom[15007] <= 10'b1000101100;
    pxcRom[15008] <= 10'b1000101100;
    pxcRom[15009] <= 10'b1000101100;
    pxcRom[15010] <= 10'b1000101100;
    pxcRom[15011] <= 10'b1000101100;
    pxcRom[15012] <= 10'b1000101100;
    pxcRom[15013] <= 10'b1000101100;
    pxcRom[15014] <= 10'b1000101100;
    pxcRom[15015] <= 10'b1000101100;
    pxcRom[15016] <= 10'b1000101100;
    pxcRom[15017] <= 10'b1000101100;
    pxcRom[15018] <= 10'b0111000101;
    pxcRom[15019] <= 10'b0110011111;
    pxcRom[15020] <= 10'b0110000011;
    pxcRom[15021] <= 10'b0101101111;
    pxcRom[15022] <= 10'b0101100011;
    pxcRom[15023] <= 10'b0101100000;
    pxcRom[15024] <= 10'b0101111010;
    pxcRom[15025] <= 10'b0110001000;
    pxcRom[15026] <= 10'b0110100111;
    pxcRom[15027] <= 10'b0111100101;
    pxcRom[15028] <= 10'b0111100101;
    pxcRom[15029] <= 10'b1000101100;
    pxcRom[15030] <= 10'b1000101100;
    pxcRom[15031] <= 10'b1000101100;
    pxcRom[15032] <= 10'b1000101100;
    pxcRom[15033] <= 10'b1000101100;
    pxcRom[15034] <= 10'b1000101100;
    pxcRom[15035] <= 10'b1000101100;
    pxcRom[15036] <= 10'b1000101100;
    pxcRom[15037] <= 10'b1000101100;
    pxcRom[15038] <= 10'b1000101100;
    pxcRom[15039] <= 10'b1000101100;
    pxcRom[15040] <= 10'b1000101100;
    pxcRom[15041] <= 10'b1000101100;
    pxcRom[15042] <= 10'b1000101100;
    pxcRom[15043] <= 10'b0111010011;
    pxcRom[15044] <= 10'b0110011000;
    pxcRom[15045] <= 10'b0101010000;
    pxcRom[15046] <= 10'b0100011010;
    pxcRom[15047] <= 10'b0011101011;
    pxcRom[15048] <= 10'b0011001101;
    pxcRom[15049] <= 10'b0010111100;
    pxcRom[15050] <= 10'b0010110101;
    pxcRom[15051] <= 10'b0010110001;
    pxcRom[15052] <= 10'b0010110111;
    pxcRom[15053] <= 10'b0011001000;
    pxcRom[15054] <= 10'b0011011111;
    pxcRom[15055] <= 10'b0011111100;
    pxcRom[15056] <= 10'b0100011111;
    pxcRom[15057] <= 10'b0101010010;
    pxcRom[15058] <= 10'b0110011000;
    pxcRom[15059] <= 10'b0111111111;
    pxcRom[15060] <= 10'b1000101100;
    pxcRom[15061] <= 10'b1000101100;
    pxcRom[15062] <= 10'b1000101100;
    pxcRom[15063] <= 10'b1000101100;
    pxcRom[15064] <= 10'b1000101100;
    pxcRom[15065] <= 10'b1000101100;
    pxcRom[15066] <= 10'b1000101100;
    pxcRom[15067] <= 10'b1000101100;
    pxcRom[15068] <= 10'b1000101100;
    pxcRom[15069] <= 10'b0111100101;
    pxcRom[15070] <= 10'b0101110110;
    pxcRom[15071] <= 10'b0101000110;
    pxcRom[15072] <= 10'b0011110100;
    pxcRom[15073] <= 10'b0010111011;
    pxcRom[15074] <= 10'b0010010001;
    pxcRom[15075] <= 10'b0001101001;
    pxcRom[15076] <= 10'b0001001010;
    pxcRom[15077] <= 10'b0000110100;
    pxcRom[15078] <= 10'b0000101000;
    pxcRom[15079] <= 10'b0000100011;
    pxcRom[15080] <= 10'b0000100110;
    pxcRom[15081] <= 10'b0000110001;
    pxcRom[15082] <= 10'b0001000101;
    pxcRom[15083] <= 10'b0001100010;
    pxcRom[15084] <= 10'b0010001010;
    pxcRom[15085] <= 10'b0010111011;
    pxcRom[15086] <= 10'b0100000111;
    pxcRom[15087] <= 10'b0101010100;
    pxcRom[15088] <= 10'b0111000101;
    pxcRom[15089] <= 10'b0111111111;
    pxcRom[15090] <= 10'b1000101100;
    pxcRom[15091] <= 10'b1000101100;
    pxcRom[15092] <= 10'b1000101100;
    pxcRom[15093] <= 10'b1000101100;
    pxcRom[15094] <= 10'b1000101100;
    pxcRom[15095] <= 10'b0111111111;
    pxcRom[15096] <= 10'b0111111111;
    pxcRom[15097] <= 10'b0101111010;
    pxcRom[15098] <= 10'b0100011011;
    pxcRom[15099] <= 10'b0011011001;
    pxcRom[15100] <= 10'b0010011101;
    pxcRom[15101] <= 10'b0001110010;
    pxcRom[15102] <= 10'b0001001001;
    pxcRom[15103] <= 10'b0000101011;
    pxcRom[15104] <= 10'b0000010111;
    pxcRom[15105] <= 10'b0000001011;
    pxcRom[15106] <= 10'b0000000110;
    pxcRom[15107] <= 10'b0000000101;
    pxcRom[15108] <= 10'b0000001000;
    pxcRom[15109] <= 10'b0000010000;
    pxcRom[15110] <= 10'b0000011111;
    pxcRom[15111] <= 10'b0000110111;
    pxcRom[15112] <= 10'b0001011010;
    pxcRom[15113] <= 10'b0010000101;
    pxcRom[15114] <= 10'b0011000011;
    pxcRom[15115] <= 10'b0100001101;
    pxcRom[15116] <= 10'b0101101001;
    pxcRom[15117] <= 10'b0111000101;
    pxcRom[15118] <= 10'b1000101100;
    pxcRom[15119] <= 10'b1000101100;
    pxcRom[15120] <= 10'b1000101100;
    pxcRom[15121] <= 10'b1000101100;
    pxcRom[15122] <= 10'b1000101100;
    pxcRom[15123] <= 10'b0111010011;
    pxcRom[15124] <= 10'b0101101100;
    pxcRom[15125] <= 10'b0100011001;
    pxcRom[15126] <= 10'b0011010101;
    pxcRom[15127] <= 10'b0010011011;
    pxcRom[15128] <= 10'b0001101001;
    pxcRom[15129] <= 10'b0001000010;
    pxcRom[15130] <= 10'b0000100011;
    pxcRom[15131] <= 10'b0000010000;
    pxcRom[15132] <= 10'b0000001001;
    pxcRom[15133] <= 10'b0000001000;
    pxcRom[15134] <= 10'b0000001001;
    pxcRom[15135] <= 10'b0000001011;
    pxcRom[15136] <= 10'b0000001011;
    pxcRom[15137] <= 10'b0000001110;
    pxcRom[15138] <= 10'b0000010110;
    pxcRom[15139] <= 10'b0000101001;
    pxcRom[15140] <= 10'b0001000101;
    pxcRom[15141] <= 10'b0001101101;
    pxcRom[15142] <= 10'b0010100011;
    pxcRom[15143] <= 10'b0011101101;
    pxcRom[15144] <= 10'b0101001100;
    pxcRom[15145] <= 10'b0110111001;
    pxcRom[15146] <= 10'b1000101100;
    pxcRom[15147] <= 10'b1000101100;
    pxcRom[15148] <= 10'b1000101100;
    pxcRom[15149] <= 10'b1000101100;
    pxcRom[15150] <= 10'b1000101100;
    pxcRom[15151] <= 10'b0110101111;
    pxcRom[15152] <= 10'b0101000000;
    pxcRom[15153] <= 10'b0011100011;
    pxcRom[15154] <= 10'b0010100110;
    pxcRom[15155] <= 10'b0001110001;
    pxcRom[15156] <= 10'b0001000101;
    pxcRom[15157] <= 10'b0000100100;
    pxcRom[15158] <= 10'b0000010010;
    pxcRom[15159] <= 10'b0000001100;
    pxcRom[15160] <= 10'b0000010000;
    pxcRom[15161] <= 10'b0000011010;
    pxcRom[15162] <= 10'b0000100101;
    pxcRom[15163] <= 10'b0000101000;
    pxcRom[15164] <= 10'b0000100000;
    pxcRom[15165] <= 10'b0000010111;
    pxcRom[15166] <= 10'b0000010110;
    pxcRom[15167] <= 10'b0000100001;
    pxcRom[15168] <= 10'b0000111100;
    pxcRom[15169] <= 10'b0001100010;
    pxcRom[15170] <= 10'b0010011001;
    pxcRom[15171] <= 10'b0011100101;
    pxcRom[15172] <= 10'b0101001000;
    pxcRom[15173] <= 10'b0110111001;
    pxcRom[15174] <= 10'b1000101100;
    pxcRom[15175] <= 10'b1000101100;
    pxcRom[15176] <= 10'b1000101100;
    pxcRom[15177] <= 10'b1000101100;
    pxcRom[15178] <= 10'b1000101100;
    pxcRom[15179] <= 10'b0101111010;
    pxcRom[15180] <= 10'b0100001010;
    pxcRom[15181] <= 10'b0010111100;
    pxcRom[15182] <= 10'b0010000110;
    pxcRom[15183] <= 10'b0001010011;
    pxcRom[15184] <= 10'b0000101110;
    pxcRom[15185] <= 10'b0000010110;
    pxcRom[15186] <= 10'b0000001110;
    pxcRom[15187] <= 10'b0000010100;
    pxcRom[15188] <= 10'b0000100111;
    pxcRom[15189] <= 10'b0001000010;
    pxcRom[15190] <= 10'b0001010110;
    pxcRom[15191] <= 10'b0001001001;
    pxcRom[15192] <= 10'b0000101110;
    pxcRom[15193] <= 10'b0000011001;
    pxcRom[15194] <= 10'b0000010011;
    pxcRom[15195] <= 10'b0000011100;
    pxcRom[15196] <= 10'b0000110110;
    pxcRom[15197] <= 10'b0001011111;
    pxcRom[15198] <= 10'b0010010111;
    pxcRom[15199] <= 10'b0011100010;
    pxcRom[15200] <= 10'b0101000110;
    pxcRom[15201] <= 10'b0110101111;
    pxcRom[15202] <= 10'b0111111111;
    pxcRom[15203] <= 10'b1000101100;
    pxcRom[15204] <= 10'b1000101100;
    pxcRom[15205] <= 10'b1000101100;
    pxcRom[15206] <= 10'b0111010011;
    pxcRom[15207] <= 10'b0101011001;
    pxcRom[15208] <= 10'b0011101011;
    pxcRom[15209] <= 10'b0010100010;
    pxcRom[15210] <= 10'b0001101101;
    pxcRom[15211] <= 10'b0001000000;
    pxcRom[15212] <= 10'b0000100000;
    pxcRom[15213] <= 10'b0000010001;
    pxcRom[15214] <= 10'b0000010011;
    pxcRom[15215] <= 10'b0000100110;
    pxcRom[15216] <= 10'b0001001010;
    pxcRom[15217] <= 10'b0001110000;
    pxcRom[15218] <= 10'b0001101101;
    pxcRom[15219] <= 10'b0001000101;
    pxcRom[15220] <= 10'b0000100100;
    pxcRom[15221] <= 10'b0000010001;
    pxcRom[15222] <= 10'b0000001101;
    pxcRom[15223] <= 10'b0000011001;
    pxcRom[15224] <= 10'b0000110110;
    pxcRom[15225] <= 10'b0001100100;
    pxcRom[15226] <= 10'b0010100000;
    pxcRom[15227] <= 10'b0011101100;
    pxcRom[15228] <= 10'b0101100000;
    pxcRom[15229] <= 10'b0111000101;
    pxcRom[15230] <= 10'b0111111111;
    pxcRom[15231] <= 10'b1000101100;
    pxcRom[15232] <= 10'b1000101100;
    pxcRom[15233] <= 10'b1000101100;
    pxcRom[15234] <= 10'b0111010011;
    pxcRom[15235] <= 10'b0100111010;
    pxcRom[15236] <= 10'b0011011000;
    pxcRom[15237] <= 10'b0010010111;
    pxcRom[15238] <= 10'b0001100000;
    pxcRom[15239] <= 10'b0000110101;
    pxcRom[15240] <= 10'b0000011011;
    pxcRom[15241] <= 10'b0000010010;
    pxcRom[15242] <= 10'b0000011011;
    pxcRom[15243] <= 10'b0000110110;
    pxcRom[15244] <= 10'b0001011010;
    pxcRom[15245] <= 10'b0001100011;
    pxcRom[15246] <= 10'b0001001001;
    pxcRom[15247] <= 10'b0000101011;
    pxcRom[15248] <= 10'b0000010100;
    pxcRom[15249] <= 10'b0000001001;
    pxcRom[15250] <= 10'b0000001011;
    pxcRom[15251] <= 10'b0000011100;
    pxcRom[15252] <= 10'b0000111101;
    pxcRom[15253] <= 10'b0001110010;
    pxcRom[15254] <= 10'b0010110010;
    pxcRom[15255] <= 10'b0100000001;
    pxcRom[15256] <= 10'b0101111010;
    pxcRom[15257] <= 10'b1000101100;
    pxcRom[15258] <= 10'b1000101100;
    pxcRom[15259] <= 10'b1000101100;
    pxcRom[15260] <= 10'b1000101100;
    pxcRom[15261] <= 10'b1000101100;
    pxcRom[15262] <= 10'b0111100101;
    pxcRom[15263] <= 10'b0100111110;
    pxcRom[15264] <= 10'b0011010000;
    pxcRom[15265] <= 10'b0010001101;
    pxcRom[15266] <= 10'b0001011011;
    pxcRom[15267] <= 10'b0000110010;
    pxcRom[15268] <= 10'b0000011010;
    pxcRom[15269] <= 10'b0000010100;
    pxcRom[15270] <= 10'b0000011110;
    pxcRom[15271] <= 10'b0000110010;
    pxcRom[15272] <= 10'b0000111101;
    pxcRom[15273] <= 10'b0000110110;
    pxcRom[15274] <= 10'b0000100110;
    pxcRom[15275] <= 10'b0000010101;
    pxcRom[15276] <= 10'b0000001001;
    pxcRom[15277] <= 10'b0000000101;
    pxcRom[15278] <= 10'b0000001100;
    pxcRom[15279] <= 10'b0000100011;
    pxcRom[15280] <= 10'b0001001110;
    pxcRom[15281] <= 10'b0010001000;
    pxcRom[15282] <= 10'b0011001001;
    pxcRom[15283] <= 10'b0100011010;
    pxcRom[15284] <= 10'b0110001000;
    pxcRom[15285] <= 10'b0111111111;
    pxcRom[15286] <= 10'b0111111111;
    pxcRom[15287] <= 10'b1000101100;
    pxcRom[15288] <= 10'b1000101100;
    pxcRom[15289] <= 10'b1000101100;
    pxcRom[15290] <= 10'b0111111111;
    pxcRom[15291] <= 10'b0101000000;
    pxcRom[15292] <= 10'b0011010011;
    pxcRom[15293] <= 10'b0010010000;
    pxcRom[15294] <= 10'b0001011111;
    pxcRom[15295] <= 10'b0000110110;
    pxcRom[15296] <= 10'b0000011110;
    pxcRom[15297] <= 10'b0000010101;
    pxcRom[15298] <= 10'b0000011001;
    pxcRom[15299] <= 10'b0000100000;
    pxcRom[15300] <= 10'b0000100000;
    pxcRom[15301] <= 10'b0000011011;
    pxcRom[15302] <= 10'b0000010100;
    pxcRom[15303] <= 10'b0000001100;
    pxcRom[15304] <= 10'b0000000101;
    pxcRom[15305] <= 10'b0000000100;
    pxcRom[15306] <= 10'b0000010001;
    pxcRom[15307] <= 10'b0000110001;
    pxcRom[15308] <= 10'b0001100100;
    pxcRom[15309] <= 10'b0010100001;
    pxcRom[15310] <= 10'b0011100100;
    pxcRom[15311] <= 10'b0100101111;
    pxcRom[15312] <= 10'b0110011111;
    pxcRom[15313] <= 10'b0111111111;
    pxcRom[15314] <= 10'b0111111111;
    pxcRom[15315] <= 10'b1000101100;
    pxcRom[15316] <= 10'b1000101100;
    pxcRom[15317] <= 10'b1000101100;
    pxcRom[15318] <= 10'b0111111111;
    pxcRom[15319] <= 10'b0101010010;
    pxcRom[15320] <= 10'b0011100000;
    pxcRom[15321] <= 10'b0010011110;
    pxcRom[15322] <= 10'b0001101011;
    pxcRom[15323] <= 10'b0001000010;
    pxcRom[15324] <= 10'b0000100111;
    pxcRom[15325] <= 10'b0000011010;
    pxcRom[15326] <= 10'b0000010111;
    pxcRom[15327] <= 10'b0000010111;
    pxcRom[15328] <= 10'b0000010111;
    pxcRom[15329] <= 10'b0000010101;
    pxcRom[15330] <= 10'b0000010010;
    pxcRom[15331] <= 10'b0000001011;
    pxcRom[15332] <= 10'b0000000101;
    pxcRom[15333] <= 10'b0000000111;
    pxcRom[15334] <= 10'b0000011001;
    pxcRom[15335] <= 10'b0001000011;
    pxcRom[15336] <= 10'b0001111010;
    pxcRom[15337] <= 10'b0010111001;
    pxcRom[15338] <= 10'b0011110101;
    pxcRom[15339] <= 10'b0100110101;
    pxcRom[15340] <= 10'b0110100111;
    pxcRom[15341] <= 10'b0111111111;
    pxcRom[15342] <= 10'b0111100101;
    pxcRom[15343] <= 10'b1000101100;
    pxcRom[15344] <= 10'b1000101100;
    pxcRom[15345] <= 10'b1000101100;
    pxcRom[15346] <= 10'b1000101100;
    pxcRom[15347] <= 10'b0101101100;
    pxcRom[15348] <= 10'b0011111010;
    pxcRom[15349] <= 10'b0010110110;
    pxcRom[15350] <= 10'b0010000100;
    pxcRom[15351] <= 10'b0001011001;
    pxcRom[15352] <= 10'b0000111010;
    pxcRom[15353] <= 10'b0000101001;
    pxcRom[15354] <= 10'b0000100001;
    pxcRom[15355] <= 10'b0000011110;
    pxcRom[15356] <= 10'b0000011110;
    pxcRom[15357] <= 10'b0000100000;
    pxcRom[15358] <= 10'b0000011001;
    pxcRom[15359] <= 10'b0000001110;
    pxcRom[15360] <= 10'b0000000111;
    pxcRom[15361] <= 10'b0000001100;
    pxcRom[15362] <= 10'b0000100110;
    pxcRom[15363] <= 10'b0001010100;
    pxcRom[15364] <= 10'b0010001111;
    pxcRom[15365] <= 10'b0011000111;
    pxcRom[15366] <= 10'b0011111101;
    pxcRom[15367] <= 10'b0101000101;
    pxcRom[15368] <= 10'b0110100111;
    pxcRom[15369] <= 10'b0111111111;
    pxcRom[15370] <= 10'b0111111111;
    pxcRom[15371] <= 10'b1000101100;
    pxcRom[15372] <= 10'b1000101100;
    pxcRom[15373] <= 10'b1000101100;
    pxcRom[15374] <= 10'b0111111111;
    pxcRom[15375] <= 10'b0110010010;
    pxcRom[15376] <= 10'b0100101010;
    pxcRom[15377] <= 10'b0011011100;
    pxcRom[15378] <= 10'b0010100111;
    pxcRom[15379] <= 10'b0001111100;
    pxcRom[15380] <= 10'b0001011101;
    pxcRom[15381] <= 10'b0001001000;
    pxcRom[15382] <= 10'b0000111101;
    pxcRom[15383] <= 10'b0000111011;
    pxcRom[15384] <= 10'b0000111001;
    pxcRom[15385] <= 10'b0000110010;
    pxcRom[15386] <= 10'b0000100000;
    pxcRom[15387] <= 10'b0000010000;
    pxcRom[15388] <= 10'b0000001011;
    pxcRom[15389] <= 10'b0000010101;
    pxcRom[15390] <= 10'b0000110100;
    pxcRom[15391] <= 10'b0001100011;
    pxcRom[15392] <= 10'b0010010110;
    pxcRom[15393] <= 10'b0011001110;
    pxcRom[15394] <= 10'b0100001111;
    pxcRom[15395] <= 10'b0101001110;
    pxcRom[15396] <= 10'b0110101111;
    pxcRom[15397] <= 10'b0111111111;
    pxcRom[15398] <= 10'b1000101100;
    pxcRom[15399] <= 10'b1000101100;
    pxcRom[15400] <= 10'b0111111111;
    pxcRom[15401] <= 10'b1000101100;
    pxcRom[15402] <= 10'b0111111111;
    pxcRom[15403] <= 10'b0111000101;
    pxcRom[15404] <= 10'b0101010110;
    pxcRom[15405] <= 10'b0100010000;
    pxcRom[15406] <= 10'b0011011001;
    pxcRom[15407] <= 10'b0010110000;
    pxcRom[15408] <= 10'b0010010000;
    pxcRom[15409] <= 10'b0001111001;
    pxcRom[15410] <= 10'b0001101011;
    pxcRom[15411] <= 10'b0001100010;
    pxcRom[15412] <= 10'b0001010101;
    pxcRom[15413] <= 10'b0000111101;
    pxcRom[15414] <= 10'b0000100011;
    pxcRom[15415] <= 10'b0000010100;
    pxcRom[15416] <= 10'b0000010010;
    pxcRom[15417] <= 10'b0000100001;
    pxcRom[15418] <= 10'b0001000001;
    pxcRom[15419] <= 10'b0001101101;
    pxcRom[15420] <= 10'b0010011101;
    pxcRom[15421] <= 10'b0011010001;
    pxcRom[15422] <= 10'b0100001000;
    pxcRom[15423] <= 10'b0101000101;
    pxcRom[15424] <= 10'b0110011111;
    pxcRom[15425] <= 10'b0111010011;
    pxcRom[15426] <= 10'b1000101100;
    pxcRom[15427] <= 10'b1000101100;
    pxcRom[15428] <= 10'b1000101100;
    pxcRom[15429] <= 10'b1000101100;
    pxcRom[15430] <= 10'b1000101100;
    pxcRom[15431] <= 10'b0111010011;
    pxcRom[15432] <= 10'b0110000011;
    pxcRom[15433] <= 10'b0101000001;
    pxcRom[15434] <= 10'b0100010000;
    pxcRom[15435] <= 10'b0011101010;
    pxcRom[15436] <= 10'b0011001011;
    pxcRom[15437] <= 10'b0010110110;
    pxcRom[15438] <= 10'b0010011100;
    pxcRom[15439] <= 10'b0010000011;
    pxcRom[15440] <= 10'b0001011111;
    pxcRom[15441] <= 10'b0000111100;
    pxcRom[15442] <= 10'b0000100100;
    pxcRom[15443] <= 10'b0000011001;
    pxcRom[15444] <= 10'b0000011011;
    pxcRom[15445] <= 10'b0000101110;
    pxcRom[15446] <= 10'b0001001011;
    pxcRom[15447] <= 10'b0001110010;
    pxcRom[15448] <= 10'b0010011101;
    pxcRom[15449] <= 10'b0011010011;
    pxcRom[15450] <= 10'b0100000110;
    pxcRom[15451] <= 10'b0101000001;
    pxcRom[15452] <= 10'b0110000011;
    pxcRom[15453] <= 10'b0111000101;
    pxcRom[15454] <= 10'b1000101100;
    pxcRom[15455] <= 10'b1000101100;
    pxcRom[15456] <= 10'b1000101100;
    pxcRom[15457] <= 10'b1000101100;
    pxcRom[15458] <= 10'b0111100101;
    pxcRom[15459] <= 10'b0111010011;
    pxcRom[15460] <= 10'b0110011000;
    pxcRom[15461] <= 10'b0101010010;
    pxcRom[15462] <= 10'b0100111110;
    pxcRom[15463] <= 10'b0100011101;
    pxcRom[15464] <= 10'b0011111011;
    pxcRom[15465] <= 10'b0011010111;
    pxcRom[15466] <= 10'b0010101100;
    pxcRom[15467] <= 10'b0001111110;
    pxcRom[15468] <= 10'b0001010100;
    pxcRom[15469] <= 10'b0000110101;
    pxcRom[15470] <= 10'b0000100101;
    pxcRom[15471] <= 10'b0000011111;
    pxcRom[15472] <= 10'b0000100110;
    pxcRom[15473] <= 10'b0000110111;
    pxcRom[15474] <= 10'b0001010010;
    pxcRom[15475] <= 10'b0001110110;
    pxcRom[15476] <= 10'b0010100000;
    pxcRom[15477] <= 10'b0011001111;
    pxcRom[15478] <= 10'b0011111111;
    pxcRom[15479] <= 10'b0100110101;
    pxcRom[15480] <= 10'b0101101100;
    pxcRom[15481] <= 10'b0110101111;
    pxcRom[15482] <= 10'b1000101100;
    pxcRom[15483] <= 10'b1000101100;
    pxcRom[15484] <= 10'b1000101100;
    pxcRom[15485] <= 10'b1000101100;
    pxcRom[15486] <= 10'b1000101100;
    pxcRom[15487] <= 10'b0111100101;
    pxcRom[15488] <= 10'b0110101111;
    pxcRom[15489] <= 10'b0101100011;
    pxcRom[15490] <= 10'b0101001010;
    pxcRom[15491] <= 10'b0100011001;
    pxcRom[15492] <= 10'b0011101111;
    pxcRom[15493] <= 10'b0010111101;
    pxcRom[15494] <= 10'b0010001111;
    pxcRom[15495] <= 10'b0001100110;
    pxcRom[15496] <= 10'b0001000110;
    pxcRom[15497] <= 10'b0000110000;
    pxcRom[15498] <= 10'b0000100111;
    pxcRom[15499] <= 10'b0000100110;
    pxcRom[15500] <= 10'b0000110000;
    pxcRom[15501] <= 10'b0000111111;
    pxcRom[15502] <= 10'b0001011000;
    pxcRom[15503] <= 10'b0001111000;
    pxcRom[15504] <= 10'b0010100001;
    pxcRom[15505] <= 10'b0011001011;
    pxcRom[15506] <= 10'b0011111101;
    pxcRom[15507] <= 10'b0100101011;
    pxcRom[15508] <= 10'b0101100000;
    pxcRom[15509] <= 10'b0111000101;
    pxcRom[15510] <= 10'b1000101100;
    pxcRom[15511] <= 10'b1000101100;
    pxcRom[15512] <= 10'b1000101100;
    pxcRom[15513] <= 10'b1000101100;
    pxcRom[15514] <= 10'b1000101100;
    pxcRom[15515] <= 10'b0111111111;
    pxcRom[15516] <= 10'b0111000101;
    pxcRom[15517] <= 10'b0110000011;
    pxcRom[15518] <= 10'b0101000000;
    pxcRom[15519] <= 10'b0100000010;
    pxcRom[15520] <= 10'b0011001010;
    pxcRom[15521] <= 10'b0010011101;
    pxcRom[15522] <= 10'b0001110100;
    pxcRom[15523] <= 10'b0001010100;
    pxcRom[15524] <= 10'b0000111100;
    pxcRom[15525] <= 10'b0000101111;
    pxcRom[15526] <= 10'b0000101011;
    pxcRom[15527] <= 10'b0000101111;
    pxcRom[15528] <= 10'b0000111000;
    pxcRom[15529] <= 10'b0001000110;
    pxcRom[15530] <= 10'b0001011011;
    pxcRom[15531] <= 10'b0001111000;
    pxcRom[15532] <= 10'b0010011111;
    pxcRom[15533] <= 10'b0011000011;
    pxcRom[15534] <= 10'b0011110001;
    pxcRom[15535] <= 10'b0100100001;
    pxcRom[15536] <= 10'b0101100000;
    pxcRom[15537] <= 10'b0111010011;
    pxcRom[15538] <= 10'b1000101100;
    pxcRom[15539] <= 10'b1000101100;
    pxcRom[15540] <= 10'b1000101100;
    pxcRom[15541] <= 10'b1000101100;
    pxcRom[15542] <= 10'b1000101100;
    pxcRom[15543] <= 10'b0111111111;
    pxcRom[15544] <= 10'b0111000101;
    pxcRom[15545] <= 10'b0101101001;
    pxcRom[15546] <= 10'b0100100011;
    pxcRom[15547] <= 10'b0011100010;
    pxcRom[15548] <= 10'b0010110000;
    pxcRom[15549] <= 10'b0010000111;
    pxcRom[15550] <= 10'b0001100010;
    pxcRom[15551] <= 10'b0001001001;
    pxcRom[15552] <= 10'b0000111001;
    pxcRom[15553] <= 10'b0000110011;
    pxcRom[15554] <= 10'b0000110011;
    pxcRom[15555] <= 10'b0000110111;
    pxcRom[15556] <= 10'b0000111111;
    pxcRom[15557] <= 10'b0001001001;
    pxcRom[15558] <= 10'b0001011110;
    pxcRom[15559] <= 10'b0001111000;
    pxcRom[15560] <= 10'b0010011001;
    pxcRom[15561] <= 10'b0011000001;
    pxcRom[15562] <= 10'b0011101010;
    pxcRom[15563] <= 10'b0100010110;
    pxcRom[15564] <= 10'b0101100000;
    pxcRom[15565] <= 10'b0111010011;
    pxcRom[15566] <= 10'b1000101100;
    pxcRom[15567] <= 10'b1000101100;
    pxcRom[15568] <= 10'b1000101100;
    pxcRom[15569] <= 10'b1000101100;
    pxcRom[15570] <= 10'b1000101100;
    pxcRom[15571] <= 10'b1000101100;
    pxcRom[15572] <= 10'b0110100111;
    pxcRom[15573] <= 10'b0101001000;
    pxcRom[15574] <= 10'b0100000111;
    pxcRom[15575] <= 10'b0011010000;
    pxcRom[15576] <= 10'b0010100001;
    pxcRom[15577] <= 10'b0001111011;
    pxcRom[15578] <= 10'b0001011100;
    pxcRom[15579] <= 10'b0001001000;
    pxcRom[15580] <= 10'b0000111100;
    pxcRom[15581] <= 10'b0000111010;
    pxcRom[15582] <= 10'b0000111100;
    pxcRom[15583] <= 10'b0001000001;
    pxcRom[15584] <= 10'b0001000111;
    pxcRom[15585] <= 10'b0001010000;
    pxcRom[15586] <= 10'b0001100010;
    pxcRom[15587] <= 10'b0001111011;
    pxcRom[15588] <= 10'b0010011001;
    pxcRom[15589] <= 10'b0010111111;
    pxcRom[15590] <= 10'b0011101111;
    pxcRom[15591] <= 10'b0100011100;
    pxcRom[15592] <= 10'b0101110011;
    pxcRom[15593] <= 10'b0111111111;
    pxcRom[15594] <= 10'b1000101100;
    pxcRom[15595] <= 10'b1000101100;
    pxcRom[15596] <= 10'b1000101100;
    pxcRom[15597] <= 10'b1000101100;
    pxcRom[15598] <= 10'b0111111111;
    pxcRom[15599] <= 10'b1000101100;
    pxcRom[15600] <= 10'b0110010010;
    pxcRom[15601] <= 10'b0101000011;
    pxcRom[15602] <= 10'b0100000010;
    pxcRom[15603] <= 10'b0011010101;
    pxcRom[15604] <= 10'b0010100110;
    pxcRom[15605] <= 10'b0010000010;
    pxcRom[15606] <= 10'b0001100101;
    pxcRom[15607] <= 10'b0001010100;
    pxcRom[15608] <= 10'b0001001011;
    pxcRom[15609] <= 10'b0001001010;
    pxcRom[15610] <= 10'b0001001110;
    pxcRom[15611] <= 10'b0001010010;
    pxcRom[15612] <= 10'b0001011001;
    pxcRom[15613] <= 10'b0001011111;
    pxcRom[15614] <= 10'b0001110001;
    pxcRom[15615] <= 10'b0010001010;
    pxcRom[15616] <= 10'b0010101001;
    pxcRom[15617] <= 10'b0011010010;
    pxcRom[15618] <= 10'b0100000001;
    pxcRom[15619] <= 10'b0100111110;
    pxcRom[15620] <= 10'b0110010010;
    pxcRom[15621] <= 10'b0111111111;
    pxcRom[15622] <= 10'b1000101100;
    pxcRom[15623] <= 10'b1000101100;
    pxcRom[15624] <= 10'b1000101100;
    pxcRom[15625] <= 10'b1000101100;
    pxcRom[15626] <= 10'b1000101100;
    pxcRom[15627] <= 10'b0111111111;
    pxcRom[15628] <= 10'b0110111001;
    pxcRom[15629] <= 10'b0101110110;
    pxcRom[15630] <= 10'b0101001010;
    pxcRom[15631] <= 10'b0100101100;
    pxcRom[15632] <= 10'b0011111000;
    pxcRom[15633] <= 10'b0011010101;
    pxcRom[15634] <= 10'b0010111001;
    pxcRom[15635] <= 10'b0010100010;
    pxcRom[15636] <= 10'b0010010111;
    pxcRom[15637] <= 10'b0010010110;
    pxcRom[15638] <= 10'b0010011000;
    pxcRom[15639] <= 10'b0010011110;
    pxcRom[15640] <= 10'b0010100101;
    pxcRom[15641] <= 10'b0010101010;
    pxcRom[15642] <= 10'b0010111011;
    pxcRom[15643] <= 10'b0011010111;
    pxcRom[15644] <= 10'b0011110100;
    pxcRom[15645] <= 10'b0100011111;
    pxcRom[15646] <= 10'b0101101100;
    pxcRom[15647] <= 10'b0110111001;
    pxcRom[15648] <= 10'b1000101100;
    pxcRom[15649] <= 10'b1000101100;
    pxcRom[15650] <= 10'b1000101100;
    pxcRom[15651] <= 10'b1000101100;
    pxcRom[15652] <= 10'b1000101100;
    pxcRom[15653] <= 10'b1000101100;
    pxcRom[15654] <= 10'b1000101100;
    pxcRom[15655] <= 10'b1000101100;
    pxcRom[15656] <= 10'b1000101100;
    pxcRom[15657] <= 10'b1000101100;
    pxcRom[15658] <= 10'b0111111111;
    pxcRom[15659] <= 10'b0111111111;
    pxcRom[15660] <= 10'b0111111111;
    pxcRom[15661] <= 10'b0111010011;
    pxcRom[15662] <= 10'b0110111001;
    pxcRom[15663] <= 10'b0110100111;
    pxcRom[15664] <= 10'b0110100111;
    pxcRom[15665] <= 10'b0110101111;
    pxcRom[15666] <= 10'b0101111010;
    pxcRom[15667] <= 10'b0110001101;
    pxcRom[15668] <= 10'b0110100111;
    pxcRom[15669] <= 10'b0110100111;
    pxcRom[15670] <= 10'b0110100111;
    pxcRom[15671] <= 10'b0110100111;
    pxcRom[15672] <= 10'b0110100111;
    pxcRom[15673] <= 10'b0111010011;
    pxcRom[15674] <= 10'b0111100101;
    pxcRom[15675] <= 10'b1000101100;
    pxcRom[15676] <= 10'b1000101100;
    pxcRom[15677] <= 10'b1000101100;
    pxcRom[15678] <= 10'b1000101100;
    pxcRom[15679] <= 10'b1000101100;

  
    end
    
    assign dout = ( ena == 0 ) ? 10'b0000_0000_00 : pxcRom[addr];
    
endmodule
